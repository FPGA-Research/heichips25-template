* NGSPICE file created from heichips25_snitch_wrapper.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_2 abstract view
.subckt sg13g2_and2_2 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_2 abstract view
.subckt sg13g2_mux2_2 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_2 abstract view
.subckt sg13g2_and4_2 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

.subckt heichips25_snitch_wrapper VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_95_840 VPWR VGND sg13g2_decap_8
XFILLER_67_520 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2699 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2612 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q_D VGND net2335 net2257
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A
+ net125 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_nor2_1
XFILLER_54_258 VPWR VGND sg13g2_decap_4
XFILLER_23_623 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2547 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2613 VPWR VGND sg13g2_a22oi_1
XFILLER_23_634 VPWR VGND sg13g2_fill_2
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2_sg13g2_inv_1_Y
+ VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B
+ VGND sg13g2_inv_1
XFILLER_50_464 VPWR VGND sg13g2_decap_8
XFILLER_10_317 VPWR VGND sg13g2_decap_4
XFILLER_10_306 VPWR VGND sg13g2_fill_2
XFILLER_22_199 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1 net2998
+ VPWR i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_a221oi_1_A1_Y
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] net584 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xfanout3209 net3210 net3209 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[355\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[355\]
+ net3121 i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_105_945 VPWR VGND sg13g2_decap_8
Xfanout2508 net2511 net2508 VPWR VGND sg13g2_buf_8
XFILLER_2_527 VPWR VGND sg13g2_fill_1
XFILLER_104_444 VPWR VGND sg13g2_fill_1
Xfanout2519 net2520 net2519 VPWR VGND sg13g2_buf_8
Xhold395 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net427 sg13g2_dlygate4sd3_1
XFILLER_77_339 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2630 net2853 net3086
+ VPWR VGND sg13g2_a22oi_1
XFILLER_93_14 VPWR VGND sg13g2_decap_8
XFILLER_86_895 VPWR VGND sg13g2_decap_8
XFILLER_85_361 VPWR VGND sg13g2_fill_2
Xhold1051 data_pdata\[28\] VPWR VGND net1083 sg13g2_dlygate4sd3_1
Xhold1040 i_snitch.i_snitch_regfile.mem\[102\] VPWR VGND net1072 sg13g2_dlygate4sd3_1
Xhold1073 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1105 sg13g2_dlygate4sd3_1
XFILLER_73_534 VPWR VGND sg13g2_fill_1
XFILLER_45_236 VPWR VGND sg13g2_decap_4
Xhold1062 i_snitch.i_snitch_regfile.mem\[368\] VPWR VGND net1094 sg13g2_dlygate4sd3_1
Xhold1084 i_snitch.i_snitch_regfile.mem\[142\] VPWR VGND net1116 sg13g2_dlygate4sd3_1
Xhold1095 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1127 sg13g2_dlygate4sd3_1
XFILLER_41_475 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2357
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR net583 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
Xrebuffer7 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_Y
+ net39 VPWR VGND sg13g2_buf_2
XFILLER_47_8 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[374\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net753 net2652 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_3_56 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2918
+ sg13g2_a221oi_1
XFILLER_95_125 VPWR VGND sg13g2_fill_1
XFILLER_83_309 VPWR VGND sg13g2_fill_1
XFILLER_49_575 VPWR VGND sg13g2_fill_1
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
XFILLER_92_843 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2393
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y net3029 sg13g2_o21ai_1
XFILLER_44_280 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2458 net2250 net2369 net1267 VPWR VGND sg13g2_a22oi_1
XFILLER_66_0 VPWR VGND sg13g2_fill_2
XFILLER_9_693 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[404\] clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_99_442 VPWR VGND sg13g2_fill_2
XFILLER_99_431 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
XFILLER_102_926 VPWR VGND sg13g2_decap_8
XFILLER_99_497 VPWR VGND sg13g2_fill_2
XFILLER_101_425 VPWR VGND sg13g2_decap_8
XFILLER_87_659 VPWR VGND sg13g2_fill_2
XFILLER_74_309 VPWR VGND sg13g2_fill_2
XFILLER_83_821 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2849 net3074 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2753 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[126\] VGND sg13g2_inv_1
XFILLER_28_726 VPWR VGND sg13g2_decap_4
XFILLER_103_35 VPWR VGND sg13g2_decap_8
XFILLER_83_865 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ net1052 VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_dfrbpq_1_Q
+ net3200 VGND VPWR net431 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_43_729 VPWR VGND sg13g2_decap_8
XFILLER_51_751 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xdata_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A VPWR data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y
+ data_pdata\[21\]_sg13g2_mux2_1_A0_X VGND sg13g2_inv_1
XFILLER_7_619 VPWR VGND sg13g2_fill_1
XFILLER_12_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2468 net2283 net2389 net1251 VPWR VGND sg13g2_a22oi_1
XFILLER_3_836 VPWR VGND sg13g2_decap_8
Xfanout3006 net3011 net3006 VPWR VGND sg13g2_buf_8
Xfanout3028 net3031 net3028 VPWR VGND sg13g2_buf_8
Xfanout3017 net3018 net3017 VPWR VGND sg13g2_buf_8
Xfanout2305 net2307 net2305 VPWR VGND sg13g2_buf_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
Xfanout3039 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y net3039 VPWR VGND sg13g2_buf_8
Xfanout2316 net2320 net2316 VPWR VGND sg13g2_buf_8
XFILLER_104_252 VPWR VGND sg13g2_decap_8
XFILLER_78_637 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[74\] net2995 VPWR VGND sg13g2_nand2_1
Xfanout2327 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2327 VPWR VGND sg13g2_buf_8
Xfanout2338 net2339 net2338 VPWR VGND sg13g2_buf_8
Xfanout2349 net2352 net2349 VPWR VGND sg13g2_buf_8
XFILLER_78_659 VPWR VGND sg13g2_decap_8
XFILLER_77_114 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_74_843 VPWR VGND sg13g2_fill_1
XFILLER_74_821 VPWR VGND sg13g2_decap_8
XFILLER_46_534 VPWR VGND sg13g2_decap_4
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_37_51 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2334
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y
+ net436 VGND sg13g2_inv_1
XFILLER_74_887 VPWR VGND sg13g2_decap_4
XFILLER_46_578 VPWR VGND sg13g2_decap_8
XFILLER_27_781 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C
+ net2747 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y
+ VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y
+ sg13g2_nor4_2
XFILLER_53_94 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[424\] clknet_leaf_74_clk sg13g2_dfrbpq_1
XFILLER_14_497 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A
+ net2706 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[213\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net1132 net2441 net2268 VPWR VGND sg13g2_a22oi_1
XFILLER_6_685 VPWR VGND sg13g2_decap_8
XFILLER_5_162 VPWR VGND sg13g2_fill_2
XFILLER_5_151 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ net2500 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X
+ net2481 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] net610 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y VGND VPWR net2759 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2 net2307 sg13g2_a21oi_1
XFILLER_69_626 VPWR VGND sg13g2_fill_1
XFILLER_97_957 VPWR VGND sg13g2_decap_8
Xfanout2850 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X
+ net2850 VPWR VGND sg13g2_buf_1
XFILLER_69_659 VPWR VGND sg13g2_fill_2
XFILLER_2_880 VPWR VGND sg13g2_decap_8
Xfanout2872 net2873 net2872 VPWR VGND sg13g2_buf_8
Xfanout2861 net2865 net2861 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[256\] VGND sg13g2_inv_1
XFILLER_49_350 VPWR VGND sg13g2_fill_1
Xfanout2894 net2896 net2894 VPWR VGND sg13g2_buf_8
Xfanout2883 net2884 net2883 VPWR VGND sg13g2_buf_8
XFILLER_92_684 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_65_887 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1
+ VPWR VGND i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[104\]
+ net2952 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2465 net2860 i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
XFILLER_21_913 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X
+ net3035 net3141 net108 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1
+ VPWR VGND sg13g2_and4_1
XFILLER_71_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_924 VPWR VGND sg13g2_fill_2
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
XFILLER_106_506 VPWR VGND sg13g2_fill_2
XFILLER_88_924 VPWR VGND sg13g2_decap_8
XFILLER_0_828 VPWR VGND sg13g2_decap_8
XFILLER_101_266 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[444\] clknet_leaf_96_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2581 VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1
+ VGND net2594 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B
+ sg13g2_o21ai_1
XFILLER_55_342 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[233\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2333 net1032 net2686 net2874 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2704 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_70_323 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2465 net2865 i_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2
+ VGND VPWR net2544 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ net2552 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X net2313 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1 VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_7_449 VPWR VGND sg13g2_fill_1
XFILLER_99_35 VPWR VGND sg13g2_decap_8
XFILLER_20_990 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR net855 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_105_561 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2577 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]
+ net3173 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_79_979 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[1\]_sg13g2_and2_1_B i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q
+ net1397 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_A VPWR VGND sg13g2_and2_1
XFILLER_94_938 VPWR VGND sg13g2_decap_8
XFILLER_19_501 VPWR VGND sg13g2_fill_1
XFILLER_93_459 VPWR VGND sg13g2_decap_4
XFILLER_58_180 VPWR VGND sg13g2_decap_4
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_545 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net470 net2403 VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[25\]_sg13g2_dfrbpq_1_Q net3238 VGND VPWR rsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[25\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_64_71 VPWR VGND sg13g2_fill_1
XFILLER_62_846 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2918
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ net47 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xhold928 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] VPWR
+ VGND net960 sg13g2_dlygate4sd3_1
Xhold917 i_snitch.i_snitch_regfile.mem\[332\] VPWR VGND net949 sg13g2_dlygate4sd3_1
XFILLER_7_983 VPWR VGND sg13g2_decap_8
XFILLER_6_471 VPWR VGND sg13g2_fill_2
Xhold906 i_snitch.i_snitch_regfile.mem\[135\] VPWR VGND net938 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ sg13g2_nand3b_1
Xhold939 i_snitch.i_snitch_regfile.mem\[158\] VPWR VGND net971 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[464\] clknet_leaf_89_clk sg13g2_dfrbpq_1
XFILLER_9_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[253\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net958 net2437 net2250 VPWR VGND sg13g2_a22oi_1
XFILLER_85_927 VPWR VGND sg13g2_decap_8
Xfanout2680 data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ net2680 VPWR VGND sg13g2_buf_8
XFILLER_97_798 VPWR VGND sg13g2_decap_8
Xfanout2691 net2692 net2691 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C
+ VGND sg13g2_inv_1
XFILLER_84_448 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[440\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[440\] net3022 VPWR VGND sg13g2_nand2_1
XFILLER_93_993 VPWR VGND sg13g2_decap_8
XFILLER_52_301 VPWR VGND sg13g2_fill_2
XFILLER_25_504 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_B2_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_B2
+ net1406 VGND sg13g2_inv_1
XFILLER_25_537 VPWR VGND sg13g2_fill_2
XFILLER_37_386 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor2_1_B
+ net2584 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_80_665 VPWR VGND sg13g2_fill_2
XFILLER_100_14 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR net633 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net104 VPWR VGND sg13g2_nand2_1
XFILLER_106_336 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1
+ VGND sg13g2_inv_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1
+ net2756 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ VPWR shift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 VGND net3172 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]
+ sg13g2_o21ai_1
Xshift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2734 shift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2
+ shift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[26\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_0_625 VPWR VGND sg13g2_decap_8
XFILLER_76_905 VPWR VGND sg13g2_fill_2
XFILLER_102_586 VPWR VGND sg13g2_fill_2
XFILLER_102_575 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2577 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_91_919 VPWR VGND sg13g2_decap_8
XFILLER_90_407 VPWR VGND sg13g2_decap_8
XFILLER_84_982 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B
+ net2596 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_43_334 VPWR VGND sg13g2_decap_8
XFILLER_16_548 VPWR VGND sg13g2_fill_2
XFILLER_43_345 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0 net3119 i_snitch.i_snitch_regfile.mem\[156\]
+ i_snitch.i_snitch_regfile.mem\[188\] i_snitch.i_snitch_regfile.mem\[220\] i_snitch.i_snitch_regfile.mem\[252\]
+ net3100 i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[484\] clknet_leaf_14_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ VPWR VGND sg13g2_a22oi_1
XFILLER_7_213 VPWR VGND sg13g2_decap_8
Xdata_pdata\[27\]_sg13g2_nand2b_1_B data_pdata\[27\]_sg13g2_nand2b_1_B_Y data_pdata\[27\]
+ VPWR VGND net3158 sg13g2_nand2b_2
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_a22oi_1_B2_Y
+ net2325 net562 net2663 net2893 VPWR VGND sg13g2_a22oi_1
XFILLER_50_62 VPWR VGND sg13g2_fill_1
XFILLER_4_920 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C VPWR
+ VGND sg13g2_nor2_1
XFILLER_106_892 VPWR VGND sg13g2_decap_8
XFILLER_4_997 VPWR VGND sg13g2_decap_8
XFILLER_61_1027 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[274\]
+ net3028 i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_a21oi_1_A1_Y net2987 sg13g2_a21oi_1
XFILLER_66_448 VPWR VGND sg13g2_fill_1
XFILLER_47_640 VPWR VGND sg13g2_fill_2
XFILLER_19_320 VPWR VGND sg13g2_fill_1
XFILLER_38_139 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net827 net2665 net3041 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xdata_pdata\[26\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net819 data_pdata\[26\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_90_952 VPWR VGND sg13g2_decap_8
XFILLER_62_632 VPWR VGND sg13g2_fill_1
XFILLER_46_161 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B VPWR VGND sg13g2_or3_1
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2868
+ net2654 VPWR VGND sg13g2_nand2_1
XFILLER_22_507 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2499 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.inst_addr_o\[19\] net2525 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_62_698 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[303\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0 net3000 i_snitch.i_snitch_regfile.mem\[275\]
+ i_snitch.i_snitch_regfile.mem\[307\] i_snitch.i_snitch_regfile.mem\[339\] i_snitch.i_snitch_regfile.mem\[371\]
+ net2976 i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_34_389 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2557 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_562 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y
+ sg13g2_o21ai_1
Xhold703 data_pdata\[1\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net735 sg13g2_dlygate4sd3_1
Xhold714 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net746 sg13g2_dlygate4sd3_1
Xhold725 i_snitch.i_snitch_regfile.mem\[439\] VPWR VGND net757 sg13g2_dlygate4sd3_1
Xhold736 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\] VPWR
+ VGND net768 sg13g2_dlygate4sd3_1
Xshift_reg_q\[22\]_sg13g2_nor2_1_A net541 net2734 shift_reg_q\[22\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xhold758 i_snitch.i_snitch_regfile.mem\[184\] VPWR VGND net790 sg13g2_dlygate4sd3_1
Xhold769 i_snitch.i_snitch_regfile.mem\[438\] VPWR VGND net801 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[95\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[95\]
+ i_snitch.i_snitch_regfile.mem\[127\] net3124 i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xhold747 i_snitch.i_snitch_regfile.mem\[425\] VPWR VGND net779 sg13g2_dlygate4sd3_1
Xcnt_q\[2\]_sg13g2_a22oi_1_B2 cnt_q\[2\]_sg13g2_a22oi_1_B2_Y cnt_q\[2\]_sg13g2_a22oi_1_B2_B1
+ net448 cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 net1 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_58_916 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[285\] net3028 VPWR VGND sg13g2_nand2_1
XFILLER_85_724 VPWR VGND sg13g2_fill_2
XFILLER_73_919 VPWR VGND sg13g2_decap_8
XFILLER_84_256 VPWR VGND sg13g2_fill_2
XFILLER_77_1012 VPWR VGND sg13g2_decap_8
XFILLER_65_492 VPWR VGND sg13g2_decap_8
XFILLER_53_621 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C_sg13g2_or4_1_X
+ net3083 net3076 net3079 net3081 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C
+ VPWR VGND sg13g2_or4_1
XFILLER_81_963 VPWR VGND sg13g2_decap_8
Xcnt_q\[2\]_sg13g2_nand3_1_A net543 net500 net448 cnt_q\[2\]_sg13g2_nand3_1_A_Y VPWR
+ VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0 net3121 i_snitch.i_snitch_regfile.mem\[394\]
+ i_snitch.i_snitch_regfile.mem\[426\] i_snitch.i_snitch_regfile.mem\[458\] i_snitch.i_snitch_regfile.mem\[490\]
+ net3110 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[18\]_sg13g2_a21oi_1_A2 VGND VPWR net3156 data_pdata\[18\] data_pdata\[18\]_sg13g2_a21oi_1_A2_Y
+ net3150 sg13g2_a21oi_1
XFILLER_106_133 VPWR VGND sg13g2_decap_8
XFILLER_20_21 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2547 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2613 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_96_14 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[428\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net936 net2692 net2863 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2886
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_0_400 VPWR VGND sg13g2_decap_8
XFILLER_1_923 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor3_1_A net1353 net2866 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_103_851 VPWR VGND sg13g2_decap_8
XFILLER_88_562 VPWR VGND sg13g2_fill_2
XFILLER_88_540 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_102_350 VPWR VGND sg13g2_decap_8
XFILLER_75_201 VPWR VGND sg13g2_fill_1
Xdata_pdata\[22\]_sg13g2_mux2_1_A1 rsp_data_q\[22\] net798 net3050 data_pdata\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_48_426 VPWR VGND sg13g2_fill_2
XFILLER_76_746 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[323\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_21_1022 VPWR VGND sg13g2_decap_8
XFILLER_75_289 VPWR VGND sg13g2_fill_2
XFILLER_17_857 VPWR VGND sg13g2_fill_2
XFILLER_72_985 VPWR VGND sg13g2_fill_2
XFILLER_72_974 VPWR VGND sg13g2_fill_1
XFILLER_71_451 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_43_164 VPWR VGND sg13g2_decap_8
XFILLER_32_849 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_nand2_2
XFILLER_84_9 VPWR VGND sg13g2_fill_1
XFILLER_61_50 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2716 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2777
+ net2662 VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[11\]_sg13g2_a22oi_1_A1 shift_reg_q\[11\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_mux2_1_A1_1_X
+ net3055 net3045 shift_reg_q\[11\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2639 i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xshift_reg_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2733 shift_reg_q\[14\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[10\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[10\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_98_359 VPWR VGND sg13g2_decap_8
XFILLER_6_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_437 VPWR VGND sg13g2_decap_8
XFILLER_39_448 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[8\] net770 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xrebuffer17 i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B net49 VPWR VGND
+ sg13g2_buf_1
Xrebuffer28 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ net60 VPWR VGND sg13g2_buf_1
Xrebuffer39 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 net71 VPWR
+ VGND sg13g2_buf_1
XFILLER_63_941 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2594 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C
+ VPWR VGND sg13g2_nor2_1
XFILLER_50_602 VPWR VGND sg13g2_fill_2
XFILLER_96_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2771
+ net2657 VPWR VGND sg13g2_nand2_1
XFILLER_22_337 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[448\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2372 net742 net2903 net2739 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2876
+ net2668 VPWR VGND sg13g2_nand2_1
Xhold511 cnt_q\[1\] VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold500 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net532 sg13g2_dlygate4sd3_1
Xhold533 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\] VPWR
+ VGND net565 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xhold544 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\] VPWR
+ VGND net576 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q net3308 VGND VPWR i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[343\] clknet_leaf_66_clk sg13g2_dfrbpq_1
Xhold522 i_snitch.i_snitch_lsu.metadata_q\[0\] VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold566 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\] VPWR
+ VGND net598 sg13g2_dlygate4sd3_1
Xhold588 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\] VPWR
+ VGND net620 sg13g2_dlygate4sd3_1
Xhold577 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] VPWR
+ VGND net609 sg13g2_dlygate4sd3_1
Xhold555 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\] VPWR
+ VGND net587 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_35 VPWR VGND sg13g2_decap_8
XFILLER_103_147 VPWR VGND sg13g2_decap_8
XFILLER_89_348 VPWR VGND sg13g2_decap_8
Xhold599 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net631 sg13g2_dlygate4sd3_1
XFILLER_98_871 VPWR VGND sg13g2_decap_8
Xhold1200 i_snitch.i_snitch_regfile.mem\[319\] VPWR VGND net1232 sg13g2_dlygate4sd3_1
XFILLER_100_854 VPWR VGND sg13g2_decap_8
Xhold1233 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\] VPWR
+ VGND net1265 sg13g2_dlygate4sd3_1
Xhold1222 i_snitch.i_snitch_regfile.mem\[288\] VPWR VGND net1254 sg13g2_dlygate4sd3_1
Xhold1211 i_snitch.i_snitch_regfile.mem\[304\] VPWR VGND net1243 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_Y
+ net2554 net2602 net2599 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nand3_1
Xhold1266 rsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1298
+ sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_57_256 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q net3251 VGND VPWR i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.gpr_waddr\[5\] clknet_leaf_15_clk sg13g2_dfrbpq_1
Xhold1255 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\] VPWR
+ VGND net1287 sg13g2_dlygate4sd3_1
Xhold1244 i_snitch.i_snitch_regfile.mem\[189\] VPWR VGND net1276 sg13g2_dlygate4sd3_1
Xhold1299 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[0\] VPWR VGND net1331 sg13g2_dlygate4sd3_1
XFILLER_57_289 VPWR VGND sg13g2_decap_8
Xhold1277 i_snitch.i_snitch_regfile.mem\[163\] VPWR VGND net1309 sg13g2_dlygate4sd3_1
Xhold1288 i_snitch.i_snitch_regfile.mem\[292\] VPWR VGND net1320 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2420 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2385
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_and2_1_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y
+ i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B VPWR VGND sg13g2_and2_2
XFILLER_13_337 VPWR VGND sg13g2_decap_8
XFILLER_13_348 VPWR VGND sg13g2_fill_2
XFILLER_15_43 VPWR VGND sg13g2_fill_2
XFILLER_25_186 VPWR VGND sg13g2_decap_4
XFILLER_40_134 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2473
+ net2263 net2668 net2798 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_114_clk clknet_5_16__leaf_clk clknet_leaf_114_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D
+ net2579 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ sg13g2_nor4_2
XFILLER_31_75 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2856
+ net2669 VPWR VGND sg13g2_nand2_1
Xstrb_out_sg13g2_inv_1_Y VPWR strb_out strb_out_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y net3008 sg13g2_o21ai_1
Xoutput20 net20 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_720 VPWR VGND sg13g2_decap_8
XFILLER_89_860 VPWR VGND sg13g2_decap_8
XFILLER_0_230 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y i_snitch.pc_d\[15\] i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2 net2308 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_49_713 VPWR VGND sg13g2_fill_2
XFILLER_0_285 VPWR VGND sg13g2_decap_8
XFILLER_1_797 VPWR VGND sg13g2_decap_8
XFILLER_63_215 VPWR VGND sg13g2_decap_8
XFILLER_17_632 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[468\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net905 net2671 net2741 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2456 VPWR VGND sg13g2_nand2_1
XFILLER_72_771 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[363\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_31_156 VPWR VGND sg13g2_fill_1
XFILLER_31_167 VPWR VGND sg13g2_fill_1
XFILLER_32_668 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net732 net2665 net2888 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_105_clk clknet_5_18__leaf_clk clknet_leaf_105_clk VPWR VGND sg13g2_buf_8
XFILLER_12_370 VPWR VGND sg13g2_fill_2
XFILLER_12_381 VPWR VGND sg13g2_fill_2
XFILLER_13_893 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2366
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2709 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_657 VPWR VGND sg13g2_fill_1
XFILLER_4_580 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[359\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[359\] net2800 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_94_351 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B
+ net2515 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_39_245 VPWR VGND sg13g2_decap_8
XFILLER_95_896 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ net1323 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2329
+ sg13g2_o21ai_1
Xdata_pdata\[29\]_sg13g2_mux2_1_A1 rsp_data_q\[29\] net846 net3049 data_pdata\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_36_974 VPWR VGND sg13g2_fill_1
Xi_snitch.inst_addr_o\[23\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[23\]
+ i_snitch.inst_addr_o\[23\] clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_50_410 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 net70 VPWR VGND
+ sg13g2_nand2_2
XFILLER_23_668 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2555 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2745 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X
+ net2928 net2924 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B
+ VPWR VGND sg13g2_and4_1
XFILLER_105_924 VPWR VGND sg13g2_decap_8
Xfanout2509 net2511 net2509 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2453 VPWR VGND sg13g2_nand2_1
XFILLER_81_1019 VPWR VGND sg13g2_decap_8
Xhold396 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\] VPWR
+ VGND net428 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[488\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net882 net2644 net2857 VPWR VGND sg13g2_a22oi_1
Xhold1030 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1062 sg13g2_dlygate4sd3_1
XFILLER_86_874 VPWR VGND sg13g2_decap_8
XFILLER_85_351 VPWR VGND sg13g2_decap_4
XFILLER_73_502 VPWR VGND sg13g2_fill_2
XFILLER_58_554 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[383\] clknet_leaf_71_clk sg13g2_dfrbpq_1
Xhold1041 i_snitch.i_snitch_regfile.mem\[349\] VPWR VGND net1073 sg13g2_dlygate4sd3_1
XFILLER_19_919 VPWR VGND sg13g2_fill_2
XFILLER_85_384 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_A1
+ net696 VGND sg13g2_inv_1
Xhold1074 i_snitch.i_snitch_regfile.mem\[214\] VPWR VGND net1106 sg13g2_dlygate4sd3_1
Xhold1085 i_snitch.i_snitch_regfile.mem\[54\] VPWR VGND net1117 sg13g2_dlygate4sd3_1
Xdata_pvalid_sg13g2_dfrbpq_1_Q net3250 VGND VPWR data_pvalid_sg13g2_dfrbpq_1_Q_D data_pvalid
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
Xhold1063 i_snitch.i_snitch_regfile.mem\[245\] VPWR VGND net1095 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_nand2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2844
+ sg13g2_a221oi_1
Xhold1052 i_snitch.i_snitch_regfile.mem\[206\] VPWR VGND net1084 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[172\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net705 net2692 net2775 VPWR VGND sg13g2_a22oi_1
Xhold1096 i_snitch.i_snitch_regfile.mem\[239\] VPWR VGND net1128 sg13g2_dlygate4sd3_1
XFILLER_60_218 VPWR VGND sg13g2_decap_4
XFILLER_42_911 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_o21ai_1_A1 net3100 VPWR i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[92\] net3126 sg13g2_o21ai_1
XFILLER_26_86 VPWR VGND sg13g2_fill_1
XFILLER_41_432 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ net2589 VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ net2545 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ net2699 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xrebuffer8 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y
+ net40 VPWR VGND sg13g2_buf_8
XFILLER_10_885 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[307\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2430 net2271 net2316 net1292 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net2603 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_1_594 VPWR VGND sg13g2_decap_8
XFILLER_77_852 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1 VPWR VGND net3103 net2823
+ i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[41\]
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1_Y net2826 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q net3278 VGND VPWR i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[202\] clknet_leaf_77_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1 VPWR
+ VGND net3091 net2929 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_Y
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2393
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_36_237 VPWR VGND sg13g2_fill_1
XFILLER_92_899 VPWR VGND sg13g2_decap_8
XFILLER_72_590 VPWR VGND sg13g2_decap_8
XFILLER_60_741 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_inv_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B
+ net3085 VPWR VGND sg13g2_inv_2
XFILLER_20_605 VPWR VGND sg13g2_fill_2
XFILLER_34_1021 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C i_snitch.inst_addr_o\[19\]
+ net2306 net62 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y VPWR VGND
+ sg13g2_nor3_1
XFILLER_102_905 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2516 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2427 sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[192\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2339 net1048 net2903 net2790 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2858
+ net2694 VPWR VGND sg13g2_nand2_1
XFILLER_87_649 VPWR VGND sg13g2_fill_1
XFILLER_86_137 VPWR VGND sg13g2_fill_2
XFILLER_101_459 VPWR VGND sg13g2_fill_2
XFILLER_83_800 VPWR VGND sg13g2_decap_8
XFILLER_68_885 VPWR VGND sg13g2_fill_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
XFILLER_103_14 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_inv_2
XFILLER_83_844 VPWR VGND sg13g2_decap_8
XFILLER_94_181 VPWR VGND sg13g2_fill_2
XFILLER_82_343 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2360 net821 net2643 net2770 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2545 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_23_465 VPWR VGND sg13g2_fill_2
XFILLER_10_115 VPWR VGND sg13g2_fill_1
XFILLER_11_616 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net963 net2472 net2285 VPWR VGND sg13g2_a22oi_1
XFILLER_10_159 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1409 net797 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1 net3023 i_snitch.i_snitch_regfile.mem\[150\]
+ i_snitch.i_snitch_regfile.mem\[182\] i_snitch.i_snitch_regfile.mem\[214\] i_snitch.i_snitch_regfile.mem\[246\]
+ net2994 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_6_119 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xnor2_1_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q net3271 VGND VPWR i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[222\] clknet_leaf_92_clk sg13g2_dfrbpq_1
Xfanout3007 net3010 net3007 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1 VPWR VGND net3112 net2822
+ i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[43\]
+ i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1_Y net2828 sg13g2_a221oi_1
XFILLER_3_815 VPWR VGND sg13g2_decap_8
Xfanout3018 net3025 net3018 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[197\]_sg13g2_nor3_1_A net1312 net2789 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net641 i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2402 net2795 i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D net2908
+ sg13g2_a221oi_1
XFILLER_104_231 VPWR VGND sg13g2_decap_8
Xfanout2306 net2307 net2306 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2760 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
Xfanout3029 net3031 net3029 VPWR VGND sg13g2_buf_8
Xfanout2317 net2319 net2317 VPWR VGND sg13g2_buf_8
XFILLER_105_798 VPWR VGND sg13g2_decap_8
Xfanout2339 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2339 VPWR VGND sg13g2_buf_8
Xfanout2328 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2328 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2453
+ net2262 net2667 net2786 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND net2601 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ sg13g2_o21ai_1
XFILLER_100_470 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1
+ net1089 net667 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y_sg13g2_xnor2_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_58_362 VPWR VGND sg13g2_fill_2
XFILLER_100_492 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y
+ net96 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ net2832 VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_33_207 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_nor2_1_Y
+ net2561 net123 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_14_454 VPWR VGND sg13g2_fill_1
XFILLER_18_1027 VPWR VGND sg13g2_fill_2
XFILLER_26_292 VPWR VGND sg13g2_decap_8
XFILLER_105_1008 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2849 net3074 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2752 sg13g2_a221oi_1
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_xnor2_1
XFILLER_10_693 VPWR VGND sg13g2_decap_4
XFILLER_6_642 VPWR VGND sg13g2_fill_2
XFILLER_5_130 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_req_arb.data_i\[44\]_sg13g2_nand3_1_A net3080 net2537 i_req_arb.data_i\[44\] i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_nand3_1
XFILLER_5_196 VPWR VGND sg13g2_fill_1
XFILLER_97_936 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1_Y
+ net2977 i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_nand2b_1_A_N_Y net3012 i_snitch.i_snitch_regfile.mem\[60\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net1011 net2455 net2247 VPWR VGND sg13g2_a22oi_1
Xfanout2851 net2853 net2851 VPWR VGND sg13g2_buf_8
Xfanout2862 net2864 net2862 VPWR VGND sg13g2_buf_8
Xfanout2840 net2841 net2840 VPWR VGND sg13g2_buf_8
Xfanout2873 net2874 net2873 VPWR VGND sg13g2_buf_8
Xfanout2895 net2896 net2895 VPWR VGND sg13g2_buf_8
Xfanout2884 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_X net2884
+ VPWR VGND sg13g2_buf_8
XFILLER_77_693 VPWR VGND sg13g2_fill_1
XFILLER_92_641 VPWR VGND sg13g2_decap_4
XFILLER_76_181 VPWR VGND sg13g2_fill_1
XFILLER_64_332 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net894 net2472 net2253 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VGND i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_18_760 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VGND net2593 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_92_696 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1 net3022 i_snitch.i_snitch_regfile.mem\[152\]
+ i_snitch.i_snitch_regfile.mem\[184\] i_snitch.i_snitch_regfile.mem\[216\] i_snitch.i_snitch_regfile.mem\[248\]
+ net2993 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2 VGND
+ VPWR net2963 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_18_793 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ net2697 net2749 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[242\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_17_292 VPWR VGND sg13g2_fill_2
XFILLER_60_593 VPWR VGND sg13g2_fill_1
XFILLER_20_413 VPWR VGND sg13g2_decap_8
XFILLER_32_262 VPWR VGND sg13g2_decap_4
XFILLER_20_446 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2347
+ sg13g2_o21ai_1
Xrsp_data_q\[6\]_sg13g2_dfrbpq_1_Q net3241 VGND VPWR rsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[6\] clknet_leaf_38_clk sg13g2_dfrbpq_2
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_Y
+ net3079 net3081 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_102_702 VPWR VGND sg13g2_decap_8
XFILLER_88_903 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ net84 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_58_18 VPWR VGND sg13g2_fill_2
XFILLER_0_807 VPWR VGND sg13g2_decap_8
XFILLER_87_446 VPWR VGND sg13g2_fill_1
Xcnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net500 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A VPWR VGND sg13g2_nand2_1
XFILLER_101_245 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.inst_addr_o\[27\] net2523 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_55_332 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_94_clk clknet_5_20__leaf_clk clknet_leaf_94_clk VPWR VGND sg13g2_buf_8
XFILLER_28_546 VPWR VGND sg13g2_decap_8
XFILLER_55_376 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\] net598 net2622
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_82_195 VPWR VGND sg13g2_decap_8
XFILLER_15_218 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ net3008 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y net2842 i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_38 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1362 net3064 net1153 VPWR VGND sg13g2_a22oi_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nand2b_1_B_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.inst_addr_o\[29\] net2523 VPWR VGND sg13g2_nand2_1
XFILLER_8_907 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR net648 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y
+ VPWR VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ sg13g2_nand4_1
XFILLER_11_468 VPWR VGND sg13g2_fill_2
XFILLER_99_14 VPWR VGND sg13g2_decap_8
XFILLER_87_1014 VPWR VGND sg13g2_decap_8
XFILLER_78_402 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[367\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net895 net2677 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_3_667 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2920
+ sg13g2_a221oi_1
XFILLER_79_958 VPWR VGND sg13g2_decap_8
XFILLER_78_435 VPWR VGND sg13g2_decap_8
XFILLER_94_917 VPWR VGND sg13g2_decap_8
XFILLER_78_468 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1 net2999 i_snitch.i_snitch_regfile.mem\[154\]
+ i_snitch.i_snitch_regfile.mem\[186\] i_snitch.i_snitch_regfile.mem\[218\] i_snitch.i_snitch_regfile.mem\[250\]
+ net2973 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A
+ sg13g2_or2_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_inv_1_A VPWR i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_inv_1_A_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A VGND sg13g2_inv_1
XFILLER_59_671 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[81\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[81\]
+ net2845 i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[262\] clknet_leaf_75_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_74_641 VPWR VGND sg13g2_decap_4
XFILLER_47_855 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_85_clk clknet_5_23__leaf_clk clknet_leaf_85_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2598 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_62_803 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y
+ net3093 VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ VGND i_snitch.sb_q\[13\] net2811 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A_Y net3019 sg13g2_o21ai_1
XFILLER_15_741 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[368\]
+ net3129 i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_a21oi_1_A1_Y net2943 sg13g2_a21oi_1
XFILLER_14_262 VPWR VGND sg13g2_decap_8
XFILLER_14_273 VPWR VGND sg13g2_fill_1
XFILLER_14_284 VPWR VGND sg13g2_fill_2
XFILLER_30_766 VPWR VGND sg13g2_fill_1
XFILLER_11_991 VPWR VGND sg13g2_fill_1
Xhold918 rsp_data_q\[16\] VPWR VGND net950 sg13g2_dlygate4sd3_1
Xhold907 i_snitch.i_snitch_regfile.mem\[87\] VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold929 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net961 sg13g2_dlygate4sd3_1
XFILLER_97_777 VPWR VGND sg13g2_fill_1
XFILLER_85_906 VPWR VGND sg13g2_decap_8
XFILLER_69_457 VPWR VGND sg13g2_fill_1
Xfanout2670 data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y
+ net2670 VPWR VGND sg13g2_buf_8
Xfanout2681 net2682 net2681 VPWR VGND sg13g2_buf_8
XFILLER_96_276 VPWR VGND sg13g2_fill_2
XFILLER_78_980 VPWR VGND sg13g2_decap_8
Xfanout2692 data_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2692 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_76_clk clknet_5_22__leaf_clk clknet_leaf_76_clk VPWR VGND sg13g2_buf_8
XFILLER_37_321 VPWR VGND sg13g2_fill_2
XFILLER_38_855 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y
+ VPWR VGND net2561 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_93_972 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q
+ net3228 VGND VPWR net440 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_53_803 VPWR VGND sg13g2_fill_1
XFILLER_92_471 VPWR VGND sg13g2_decap_8
XFILLER_80_622 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y net645
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 VPWR VGND sg13g2_inv_4
XFILLER_61_880 VPWR VGND sg13g2_decap_8
XFILLER_52_379 VPWR VGND sg13g2_fill_1
Xstate_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_B1 VGND VPWR net1 i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y
+ target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_106_315 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q clknet_leaf_46_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1 net3004 i_snitch.i_snitch_regfile.mem\[156\]
+ i_snitch.i_snitch_regfile.mem\[188\] i_snitch.i_snitch_regfile.mem\[220\] i_snitch.i_snitch_regfile.mem\[252\]
+ net2978 i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2 i_snitch.inst_addr_o\[15\] i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_69_39 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q net3208 VGND VPWR i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[282\] clknet_leaf_117_clk sg13g2_dfrbpq_1
XFILLER_0_604 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1 VPWR VGND net3109 net2822
+ i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[49\]
+ i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1_Y net2830 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_88_788 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_67_clk clknet_5_30__leaf_clk clknet_leaf_67_clk VPWR VGND sg13g2_buf_8
XFILLER_84_961 VPWR VGND sg13g2_decap_8
XFILLER_71_600 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[3\]_sg13g2_nor2_1_A net521 net2732 shift_reg_q\[3\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[121\]
+ net2998 i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_70_154 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_nor2_1_B i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A i_snitch.pc_d\[5\]
+ i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[417\] clknet_leaf_103_clk sg13g2_dfrbpq_1
XFILLER_43_379 VPWR VGND sg13g2_fill_2
XFILLER_24_571 VPWR VGND sg13g2_fill_2
XFILLER_34_42 VPWR VGND sg13g2_fill_1
XFILLER_34_64 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[206\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net1084 net2688 net2792 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[101\] clknet_leaf_112_clk sg13g2_dfrbpq_1
XFILLER_106_871 VPWR VGND sg13g2_decap_8
XFILLER_4_976 VPWR VGND sg13g2_decap_8
XFILLER_3_486 VPWR VGND sg13g2_fill_2
XFILLER_105_392 VPWR VGND sg13g2_decap_8
XFILLER_78_254 VPWR VGND sg13g2_fill_1
XFILLER_93_213 VPWR VGND sg13g2_fill_2
XFILLER_79_788 VPWR VGND sg13g2_decap_4
XFILLER_78_287 VPWR VGND sg13g2_fill_2
XFILLER_22_8 VPWR VGND sg13g2_fill_1
XFILLER_39_619 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ net88 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_82_909 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_58_clk clknet_5_30__leaf_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
Xdata_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 net2682 VPWR
+ data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y
+ net3068 sg13g2_o21ai_1
XFILLER_81_419 VPWR VGND sg13g2_decap_8
XFILLER_75_71 VPWR VGND sg13g2_fill_2
XFILLER_47_663 VPWR VGND sg13g2_fill_1
XFILLER_47_652 VPWR VGND sg13g2_fill_2
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_35_814 VPWR VGND sg13g2_fill_1
XFILLER_90_931 VPWR VGND sg13g2_decap_8
XFILLER_75_994 VPWR VGND sg13g2_fill_2
XFILLER_74_471 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ net2852 net3019 sg13g2_a21oi_2
XFILLER_62_622 VPWR VGND sg13g2_decap_4
XFILLER_35_836 VPWR VGND sg13g2_decap_4
XFILLER_50_839 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1 net3012 i_snitch.i_snitch_regfile.mem\[158\]
+ i_snitch.i_snitch_regfile.mem\[190\] i_snitch.i_snitch_regfile.mem\[222\] i_snitch.i_snitch_regfile.mem\[254\]
+ net2985 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_req_register.data_o\[42\]_sg13g2_mux2_1_X i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\] net3166 i_req_register.data_o\[42\]
+ VPWR VGND sg13g2_mux2_1
Xshift_reg_q\[8\]_sg13g2_dfrbpq_1_Q net3229 VGND VPWR net504 shift_reg_q\[8\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
Xhold715 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\] VPWR
+ VGND net747 sg13g2_dlygate4sd3_1
Xhold726 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] VPWR
+ VGND net758 sg13g2_dlygate4sd3_1
Xhold737 i_snitch.i_snitch_regfile.mem\[86\] VPWR VGND net769 sg13g2_dlygate4sd3_1
Xhold704 i_snitch.i_snitch_regfile.mem\[105\] VPWR VGND net736 sg13g2_dlygate4sd3_1
XFILLER_89_519 VPWR VGND sg13g2_fill_2
Xhold759 i_snitch.i_snitch_regfile.mem\[215\] VPWR VGND net791 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold748 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y VPWR VGND net780 sg13g2_dlygate4sd3_1
XFILLER_103_329 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2499 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2479 VPWR VGND sg13g2_a22oi_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
XFILLER_97_541 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2417 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xfanout3190 net3193 net3190 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[298\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[298\] net2812 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[437\] clknet_leaf_114_clk sg13g2_dfrbpq_1
XFILLER_66_950 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_49_clk clknet_5_13__leaf_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
XFILLER_38_630 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[2\]
+ VGND net2292 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_81_942 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B
+ net2719 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D_X
+ VPWR VGND sg13g2_or4_1
XFILLER_65_471 VPWR VGND sg13g2_decap_8
XFILLER_26_836 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q net3215 VGND VPWR i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[121\] clknet_leaf_112_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_80_496 VPWR VGND sg13g2_fill_2
XFILLER_52_198 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1183 net3066 rsp_data_q\[4\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y_sg13g2_nand4_1_D i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B_X
+ i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_D VPWR VGND i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y
+ sg13g2_nand4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_nand2_1_A_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_A2 net2621 sg13g2_o21ai_1
XFILLER_101_1022 VPWR VGND sg13g2_decap_8
Xi_req_arb.data_i\[40\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.pc_d\[5\] i_req_arb.data_i\[40\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
XFILLER_106_112 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_fill_1
XFILLER_84_1028 VPWR VGND sg13g2_fill_1
XFILLER_84_1017 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[20\]_sg13g2_dfrbpq_1_Q net3229 VGND VPWR net497 shift_reg_q\[20\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_1_902 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2855 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2
+ net2505 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_106_189 VPWR VGND sg13g2_decap_8
Xdata_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[2\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y data_pdata\[18\]_sg13g2_mux2_1_A0_X
+ net3150 sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_X
+ net3094 net2930 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_103_830 VPWR VGND sg13g2_decap_8
XFILLER_49_906 VPWR VGND sg13g2_fill_2
XFILLER_1_979 VPWR VGND sg13g2_decap_8
XFILLER_88_585 VPWR VGND sg13g2_decap_8
XFILLER_48_405 VPWR VGND sg13g2_decap_8
XFILLER_75_246 VPWR VGND sg13g2_fill_1
XFILLER_29_630 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2577 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xrsp_data_q\[18\]_sg13g2_dfrbpq_1_Q net3231 VGND VPWR rsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[18\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_63_419 VPWR VGND sg13g2_decap_8
XFILLER_44_622 VPWR VGND sg13g2_fill_2
XFILLER_16_313 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_nor2_1_Y i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A VPWR VGND sg13g2_nor2_2
XFILLER_43_154 VPWR VGND sg13g2_fill_1
XFILLER_16_379 VPWR VGND sg13g2_fill_1
XFILLER_101_91 VPWR VGND sg13g2_decap_8
XFILLER_8_512 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[3\] net1139 net2916 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[332\] net2952 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[457\] clknet_leaf_72_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2531 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ net2480 VPWR VGND sg13g2_a22oi_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_99_839 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[246\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net903 net2651 net2875 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[403\]
+ i_snitch.i_snitch_regfile.mem\[435\] i_snitch.i_snitch_regfile.mem\[467\] i_snitch.i_snitch_regfile.mem\[499\]
+ net3098 i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_106_690 VPWR VGND sg13g2_fill_1
XFILLER_79_552 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[69\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2408 i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nor3_1_A_Y net2451 net2782 i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_dfrbpq_1_Q_D
+ net2906 sg13g2_a221oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2700 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_94_500 VPWR VGND sg13g2_fill_1
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_94_533 VPWR VGND sg13g2_fill_1
XFILLER_67_769 VPWR VGND sg13g2_fill_2
XFILLER_67_747 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[141\] clknet_leaf_85_clk sg13g2_dfrbpq_1
Xrebuffer18 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ net50 VPWR VGND sg13g2_buf_1
XFILLER_48_950 VPWR VGND sg13g2_fill_2
Xrebuffer29 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ net61 VPWR VGND sg13g2_buf_1
XFILLER_82_739 VPWR VGND sg13g2_fill_2
XFILLER_63_931 VPWR VGND sg13g2_fill_1
XFILLER_47_482 VPWR VGND sg13g2_decap_8
XFILLER_19_173 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_62_441 VPWR VGND sg13g2_fill_2
XFILLER_47_493 VPWR VGND sg13g2_fill_1
XFILLER_34_121 VPWR VGND sg13g2_fill_1
XFILLER_62_485 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2559 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net47 net2709 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND
+ sg13g2_inv_1
Xhold501 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\] VPWR
+ VGND net533 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xhold545 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\] VPWR
+ VGND net577 sg13g2_dlygate4sd3_1
Xhold523 i_snitch.sb_q\[12\] VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold534 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\] VPWR
+ VGND net566 sg13g2_dlygate4sd3_1
Xhold512 i_snitch.sb_q\[7\] VPWR VGND net544 sg13g2_dlygate4sd3_1
XFILLER_104_627 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold578 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\] VPWR
+ VGND net610 sg13g2_dlygate4sd3_1
Xhold567 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net599 sg13g2_dlygate4sd3_1
Xhold556 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net588 sg13g2_dlygate4sd3_1
XFILLER_106_14 VPWR VGND sg13g2_decap_8
XFILLER_103_126 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VGND net2584 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_98_850 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B
+ sg13g2_nand3b_1
Xhold589 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net621 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_A1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B
+ sg13g2_a21oi_1
XFILLER_100_833 VPWR VGND sg13g2_decap_8
XFILLER_97_382 VPWR VGND sg13g2_fill_1
XFILLER_57_235 VPWR VGND sg13g2_fill_1
Xhold1201 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] VPWR
+ VGND net1233 sg13g2_dlygate4sd3_1
Xhold1234 i_snitch.i_snitch_regfile.mem\[305\] VPWR VGND net1266 sg13g2_dlygate4sd3_1
Xhold1223 i_snitch.i_snitch_regfile.mem\[435\] VPWR VGND net1255 sg13g2_dlygate4sd3_1
Xhold1212 i_snitch.i_snitch_regfile.mem\[190\] VPWR VGND net1244 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold1267 rsp_data_q\[7\] VPWR VGND net1299 sg13g2_dlygate4sd3_1
Xhold1245 i_snitch.i_snitch_regfile.mem\[483\] VPWR VGND net1277 sg13g2_dlygate4sd3_1
Xhold1256 i_snitch.i_snitch_regfile.mem\[69\] VPWR VGND net1288 sg13g2_dlygate4sd3_1
Xi_req_register.data_o\[5\]_sg13g2_mux2_1_X i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\] net3164 i_req_register.data_o\[5\]
+ VPWR VGND sg13g2_mux2_1
XFILLER_85_588 VPWR VGND sg13g2_decap_4
XFILLER_72_227 VPWR VGND sg13g2_decap_8
Xhold1278 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] VPWR
+ VGND net1310 sg13g2_dlygate4sd3_1
Xhold1289 i_snitch.i_snitch_regfile.mem\[453\] VPWR VGND net1321 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] net3174
+ sg13g2_o21ai_1
XFILLER_54_964 VPWR VGND sg13g2_fill_2
XFILLER_81_794 VPWR VGND sg13g2_fill_2
XFILLER_15_22 VPWR VGND sg13g2_fill_2
XFILLER_25_143 VPWR VGND sg13g2_decap_8
XFILLER_26_677 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[477\] clknet_leaf_96_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net1020 net2434 net2283 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2392
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2867
+ net2658 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[161\] clknet_leaf_103_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y
+ VPWR VGND net3072 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ net95 net2719 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N
+ i_snitch.consec_pc\[0\] sg13g2_a221oi_1
Xoutput21 net21 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput10 net10 uio_out[1] VPWR VGND sg13g2_buf_1
XFILLER_103_671 VPWR VGND sg13g2_fill_2
XFILLER_0_242 VPWR VGND sg13g2_decap_8
XFILLER_1_776 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2261
+ sg13g2_o21ai_1
XFILLER_56_40 VPWR VGND sg13g2_fill_2
XFILLER_36_408 VPWR VGND sg13g2_fill_2
Xdata_pdata\[19\]_sg13g2_dfrbpq_1_Q net3202 VGND VPWR net755 data_pdata\[19\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_91_569 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2 i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_B1 VPWR
+ i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_Y VGND i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_A1
+ i_snitch.pc_d\[6\] sg13g2_o21ai_1
XFILLER_56_290 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A
+ net2546 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2500 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_463 VPWR VGND sg13g2_fill_2
XFILLER_17_666 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[9\]
+ VGND net2292 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_72_794 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1349 net3063 rsp_data_q\[13\] VPWR VGND sg13g2_a22oi_1
XFILLER_13_850 VPWR VGND sg13g2_fill_1
XFILLER_13_872 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2422 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y i_snitch.pc_d\[8\] i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2 net2305 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_28_1018 VPWR VGND sg13g2_decap_8
XFILLER_97_91 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1354 net2494 net1376 VPWR VGND sg13g2_a22oi_1
XFILLER_95_875 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2321
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[68\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[68\]
+ i_snitch.i_snitch_regfile.mem\[100\] net3123 i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[497\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_94_396 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2885
+ net2659 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_a22oi_1_B2_Y
+ net2327 net671 net2434 net2245 VPWR VGND sg13g2_a22oi_1
XFILLER_51_923 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_36_997 VPWR VGND sg13g2_decap_8
XFILLER_74_1027 VPWR VGND sg13g2_fill_2
XFILLER_50_422 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[181\] clknet_leaf_98_clk sg13g2_dfrbpq_1
XFILLER_51_967 VPWR VGND sg13g2_decap_8
XFILLER_105_903 VPWR VGND sg13g2_decap_8
XFILLER_104_413 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[339\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[339\] net2947 VPWR VGND sg13g2_nand2_1
Xhold397 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net429 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_nor2_1_B
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[316\] clknet_leaf_101_clk sg13g2_dfrbpq_1
XFILLER_86_853 VPWR VGND sg13g2_decap_8
XFILLER_85_341 VPWR VGND sg13g2_fill_2
Xhold1020 rsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1052
+ sg13g2_dlygate4sd3_1
Xhold1031 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]
+ VPWR VGND net1063 sg13g2_dlygate4sd3_1
Xhold1042 i_req_arb.data_i\[44\] VPWR VGND net1074 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[105\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2410 net736 net2685 net2869 VPWR VGND sg13g2_a22oi_1
Xhold1075 rsp_data_q\[31\] VPWR VGND net1107 sg13g2_dlygate4sd3_1
XFILLER_45_216 VPWR VGND sg13g2_decap_4
Xhold1064 i_snitch.i_snitch_regfile.mem\[462\] VPWR VGND net1096 sg13g2_dlygate4sd3_1
XFILLER_93_49 VPWR VGND sg13g2_fill_2
Xhold1086 i_snitch.i_snitch_regfile.mem\[280\] VPWR VGND net1118 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net467 net2394 VPWR VGND sg13g2_nand2_1
Xhold1097 i_snitch.i_snitch_regfile.mem\[412\] VPWR VGND net1129 sg13g2_dlygate4sd3_1
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y
+ net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\] VPWR
+ VGND sg13g2_nand2_1
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VGND net75 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A
+ sg13g2_o21ai_1
XFILLER_9_128 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xrebuffer9 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1_Y
+ net41 VPWR VGND sg13g2_buf_8
Xi_snitch.inst_addr_o\[1\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.pc_d\[1\]
+ i_snitch.inst_addr_o\[1\] clknet_leaf_47_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2771
+ net2661 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2
+ VGND sg13g2_inv_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C i_snitch.inst_addr_o\[10\]
+ net2306 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2413
+ sg13g2_o21ai_1
XFILLER_69_809 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[458\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net513 net2374 VPWR VGND sg13g2_nand2_1
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_104_991 VPWR VGND sg13g2_decap_8
XFILLER_89_691 VPWR VGND sg13g2_fill_1
XFILLER_77_831 VPWR VGND sg13g2_decap_4
XFILLER_1_573 VPWR VGND sg13g2_decap_8
XFILLER_67_72 VPWR VGND sg13g2_decap_4
XFILLER_97_1027 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2478 i_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2436 net2873 i_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
XFILLER_37_717 VPWR VGND sg13g2_decap_4
XFILLER_92_878 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2431
+ net2513 VPWR VGND sg13g2_nand2_1
XFILLER_72_580 VPWR VGND sg13g2_fill_2
XFILLER_80_4 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y VPWR
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\] clknet_leaf_46_clk
+ sg13g2_dfrbpq_1
XFILLER_66_2 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q net3286 VGND VPWR i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[336\] clknet_leaf_93_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2418 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2450 net2251 net2410 net1180 VPWR VGND sg13g2_a22oi_1
XFILLER_99_444 VPWR VGND sg13g2_fill_1
XFILLER_99_433 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2490 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_inv_1_A
+ VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B
+ VGND sg13g2_inv_1
XFILLER_86_105 VPWR VGND sg13g2_fill_2
XFILLER_68_820 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B
+ net2500 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_650 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[24\]_sg13g2_a22oi_1_A1 shift_reg_q\[24\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3047 shift_reg_q\[24\] VPWR VGND sg13g2_a22oi_1
XFILLER_27_227 VPWR VGND sg13g2_fill_2
XFILLER_70_528 VPWR VGND sg13g2_decap_8
XFILLER_55_569 VPWR VGND sg13g2_decap_4
XFILLER_42_219 VPWR VGND sg13g2_decap_4
XFILLER_36_783 VPWR VGND sg13g2_fill_2
XFILLER_50_285 VPWR VGND sg13g2_decap_8
XFILLER_50_296 VPWR VGND sg13g2_fill_2
Xfanout3019 net3024 net3019 VPWR VGND sg13g2_buf_8
Xfanout3008 net3009 net3008 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1388 net2491 net1283 VPWR VGND sg13g2_a22oi_1
XFILLER_104_210 VPWR VGND sg13g2_decap_8
Xfanout2307 net106 net2307 VPWR VGND sg13g2_buf_8
XFILLER_2_348 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_105_777 VPWR VGND sg13g2_decap_8
XFILLER_78_606 VPWR VGND sg13g2_fill_2
Xfanout2318 net2319 net2318 VPWR VGND sg13g2_buf_8
Xfanout2329 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2329 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2878
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_104_287 VPWR VGND sg13g2_decap_8
XFILLER_19_706 VPWR VGND sg13g2_fill_2
XFILLER_101_994 VPWR VGND sg13g2_decap_8
XFILLER_73_311 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_X
+ net3094 net2929 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2b_1_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[356\] clknet_leaf_107_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2742
+ net2653 VPWR VGND sg13g2_nand2_1
XFILLER_14_433 VPWR VGND sg13g2_decap_8
XFILLER_42_764 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2334
+ sg13g2_o21ai_1
XFILLER_53_96 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2352 net767 net2663 net2890 VPWR VGND sg13g2_a22oi_1
XFILLER_41_263 VPWR VGND sg13g2_fill_2
Xrsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1322 net3066 rsp_data_q\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_6_676 VPWR VGND sg13g2_decap_4
XFILLER_97_915 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y net2308 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2 VPWR VGND sg13g2_nor2_1
Xfanout2830 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_A2 net2830 VPWR
+ VGND sg13g2_buf_8
Xfanout2852 net2853 net2852 VPWR VGND sg13g2_buf_2
Xfanout2863 net2864 net2863 VPWR VGND sg13g2_buf_8
Xfanout2841 net2842 net2841 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_84_609 VPWR VGND sg13g2_decap_4
Xfanout2885 net2886 net2885 VPWR VGND sg13g2_buf_8
Xfanout2896 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_X net2896
+ VPWR VGND sg13g2_buf_8
Xfanout2874 net2877 net2874 VPWR VGND sg13g2_buf_8
XFILLER_92_664 VPWR VGND sg13g2_fill_1
Xi_snitch.inst_addr_o\[16\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[16\]
+ i_snitch.inst_addr_o\[16\] clknet_leaf_57_clk sg13g2_dfrbpq_2
XFILLER_17_260 VPWR VGND sg13g2_decap_4
XFILLER_17_271 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2549 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_32_230 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2340
+ sg13g2_o21ai_1
XFILLER_71_0 VPWR VGND sg13g2_fill_2
XFILLER_99_252 VPWR VGND sg13g2_decap_8
XFILLER_99_241 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q
+ net3240 VGND VPWR net999 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3085 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2849 net3075 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2751 sg13g2_a221oi_1
XFILLER_88_959 VPWR VGND sg13g2_decap_8
XFILLER_102_758 VPWR VGND sg13g2_fill_2
XFILLER_101_224 VPWR VGND sg13g2_decap_8
XFILLER_59_138 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[376\] clknet_leaf_70_clk sg13g2_dfrbpq_2
XFILLER_96_992 VPWR VGND sg13g2_decap_8
XFILLER_28_503 VPWR VGND sg13g2_decap_8
XFILLER_95_480 VPWR VGND sg13g2_decap_4
XFILLER_68_694 VPWR VGND sg13g2_fill_1
XFILLER_67_193 VPWR VGND sg13g2_fill_2
XFILLER_56_845 VPWR VGND sg13g2_decap_4
XFILLER_83_664 VPWR VGND sg13g2_fill_2
XFILLER_55_355 VPWR VGND sg13g2_fill_2
XFILLER_70_314 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_o21ai_1_A1 net3100 VPWR i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[85\] net3120 sg13g2_o21ai_1
XFILLER_90_28 VPWR VGND sg13g2_decap_8
XFILLER_70_358 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ VGND net2717 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_23_33 VPWR VGND sg13g2_fill_2
XFILLER_23_55 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_3_646 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_79_937 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1_sg13g2_o21ai_1_Y
+ net2527 VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1
+ VGND i_snitch.inst_addr_o\[15\] i_snitch.inst_addr_o\[16\] sg13g2_o21ai_1
XFILLER_78_425 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y
+ net1253 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C
+ VPWR VGND sg13g2_nor2_1
XFILLER_65_119 VPWR VGND sg13g2_fill_1
XFILLER_101_791 VPWR VGND sg13g2_decap_8
XFILLER_94_1008 VPWR VGND sg13g2_decap_8
XFILLER_104_91 VPWR VGND sg13g2_decap_8
XFILLER_74_697 VPWR VGND sg13g2_decap_4
XFILLER_62_848 VPWR VGND sg13g2_fill_1
XFILLER_15_720 VPWR VGND sg13g2_fill_2
XFILLER_34_539 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2551 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ sg13g2_a21oi_1
XFILLER_15_731 VPWR VGND sg13g2_fill_2
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_42_572 VPWR VGND sg13g2_fill_1
Xstrb_reg_q\[1\]_sg13g2_nor2_1_A net525 net2727 strb_reg_q\[1\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C i_snitch.inst_addr_o\[1\] net2301
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
Xhold919 rsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net951 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[396\] clknet_leaf_68_clk sg13g2_dfrbpq_1
XFILLER_10_491 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q
+ net3192 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
Xhold908 i_snitch.i_snitch_regfile.mem\[270\] VPWR VGND net940 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ net2539 sg13g2_a21oi_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[185\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2442 net2266 net2342 net1188 VPWR VGND sg13g2_a22oi_1
Xshift_reg_q\[17\]_sg13g2_nor2_1_A net481 net2729 shift_reg_q\[17\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_69_414 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[340\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_97_756 VPWR VGND sg13g2_fill_2
XFILLER_96_233 VPWR VGND sg13g2_fill_2
XFILLER_96_222 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]
+ net3181 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xfanout2671 net2672 net2671 VPWR VGND sg13g2_buf_8
Xfanout2660 data_pdata\[26\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2660 VPWR
+ VGND sg13g2_buf_8
Xfanout2682 net2683 net2682 VPWR VGND sg13g2_buf_2
Xfanout2693 net2694 net2693 VPWR VGND sg13g2_buf_8
XFILLER_38_801 VPWR VGND sg13g2_fill_2
XFILLER_93_951 VPWR VGND sg13g2_decap_8
XFILLER_77_480 VPWR VGND sg13g2_fill_1
XFILLER_65_642 VPWR VGND sg13g2_fill_1
XFILLER_64_141 VPWR VGND sg13g2_fill_1
XFILLER_64_130 VPWR VGND sg13g2_decap_8
XFILLER_52_303 VPWR VGND sg13g2_fill_1
XFILLER_25_539 VPWR VGND sg13g2_fill_1
XFILLER_37_388 VPWR VGND sg13g2_fill_1
XFILLER_52_347 VPWR VGND sg13g2_fill_1
XFILLER_100_49 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1153 net3064 rsp_data_q\[11\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[215\] clknet_leaf_57_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y net3019 sg13g2_o21ai_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2594 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_88_734 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_88_778 VPWR VGND sg13g2_fill_1
XFILLER_87_277 VPWR VGND sg13g2_decap_8
XFILLER_84_940 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[4\]_sg13g2_a21oi_1_A1 VGND VPWR strb_reg_q\[4\] net3043 strb_reg_q\[4\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[4\]_sg13g2_a21oi_1_A1_B1 sg13g2_a21oi_1
XFILLER_18_33 VPWR VGND sg13g2_decap_8
XFILLER_56_664 VPWR VGND sg13g2_fill_2
XFILLER_56_653 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2737 shift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2
+ shift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[27\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_29_889 VPWR VGND sg13g2_fill_2
XFILLER_16_528 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[417\]_sg13g2_a221oi_1_A1 VPWR VGND i_snitch.i_snitch_regfile.mem\[385\]
+ net2936 net2920 i_snitch.i_snitch_regfile.mem\[417\] i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_a221oi_1_A1_Y
+ net2825 sg13g2_a221oi_1
XFILLER_55_196 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_756 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2371 net842 net2645 net2856 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1
+ net1061 net565 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2_sg13g2_a21o_1_X
+ net2536 net3086 i_req_arb.data_i\[41\] i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[470\] VGND sg13g2_inv_1
XFILLER_50_86 VPWR VGND sg13g2_fill_1
XFILLER_106_850 VPWR VGND sg13g2_decap_8
XFILLER_4_955 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net867 net2455 net2269 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1_Y
+ net2978 i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_nand2b_1_A_N_Y net3004 i_snitch.i_snitch_regfile.mem\[53\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_105_371 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_59_84 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ net1366 VGND sg13g2_inv_1
XFILLER_75_984 VPWR VGND sg13g2_fill_1
XFILLER_47_642 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ net2590 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_910 VPWR VGND sg13g2_decap_8
Xdata_pdata\[12\]_sg13g2_nor2b_1_A data_pdata\[12\] net3161 data_pdata\[12\]_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.sb_q\[8\] VGND sg13g2_inv_1
XFILLER_46_185 VPWR VGND sg13g2_decap_8
XFILLER_46_152 VPWR VGND sg13g2_decap_8
XFILLER_19_377 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[235\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_90_987 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_7_760 VPWR VGND sg13g2_decap_8
Xhold716 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net748 sg13g2_dlygate4sd3_1
Xhold727 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net759 sg13g2_dlygate4sd3_1
Xhold705 i_snitch.i_snitch_regfile.mem\[360\] VPWR VGND net737 sg13g2_dlygate4sd3_1
XFILLER_104_809 VPWR VGND sg13g2_decap_8
Xhold738 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] VPWR
+ VGND net770 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2939 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xhold749 i_snitch.i_snitch_regfile.mem\[345\] VPWR VGND net781 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_103_308 VPWR VGND sg13g2_decap_8
XFILLER_69_200 VPWR VGND sg13g2_fill_1
Xfanout3180 net3180 net3181 VPWR VGND sg13g2_buf_16
Xfanout3191 net3193 net3191 VPWR VGND sg13g2_buf_8
XFILLER_97_586 VPWR VGND sg13g2_decap_8
XFILLER_97_564 VPWR VGND sg13g2_fill_2
XFILLER_85_726 VPWR VGND sg13g2_fill_1
XFILLER_84_203 VPWR VGND sg13g2_fill_1
Xfanout2490 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y
+ net2490 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1
+ net1390 VGND sg13g2_inv_1
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_26_815 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_81_921 VPWR VGND sg13g2_decap_8
XFILLER_53_623 VPWR VGND sg13g2_fill_1
XFILLER_1_91 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_686 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2700 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D_sg13g2_a221oi_1_Y
+ VPWR VGND net2925 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B_Y
+ net2922 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ sg13g2_a221oi_1
XFILLER_53_645 VPWR VGND sg13g2_fill_1
XFILLER_52_133 VPWR VGND sg13g2_decap_4
XFILLER_38_1009 VPWR VGND sg13g2_decap_8
XFILLER_81_998 VPWR VGND sg13g2_decap_8
XFILLER_80_464 VPWR VGND sg13g2_decap_4
XFILLER_53_678 VPWR VGND sg13g2_decap_8
XFILLER_34_870 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2795 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2
+ net2506 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[73\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2354 net794 net2686 net2785 VPWR VGND sg13g2_a22oi_1
XFILLER_101_1001 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_106_168 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2594 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_96_49 VPWR VGND sg13g2_decap_8
XFILLER_1_958 VPWR VGND sg13g2_decap_8
XFILLER_103_886 VPWR VGND sg13g2_decap_8
XFILLER_88_575 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q net3305 VGND VPWR i_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[255\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_0_468 VPWR VGND sg13g2_decap_8
XFILLER_102_385 VPWR VGND sg13g2_decap_8
XFILLER_48_428 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2587 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_57_962 VPWR VGND sg13g2_fill_1
XFILLER_84_792 VPWR VGND sg13g2_fill_1
XFILLER_17_848 VPWR VGND sg13g2_fill_2
XFILLER_29_697 VPWR VGND sg13g2_decap_8
XFILLER_44_645 VPWR VGND sg13g2_fill_1
XFILLER_17_859 VPWR VGND sg13g2_fill_1
XFILLER_71_486 VPWR VGND sg13g2_decap_4
XFILLER_101_70 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2 i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y i_snitch.pc_d\[30\]
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1 i_snitch.pc_d\[24\] i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2681 data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_8_568 VPWR VGND sg13g2_decap_4
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_99_818 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2544 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_4_741 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ net2705 sg13g2_or2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B
+ net3144 net3141 VPWR VGND sg13g2_nand2_2
XFILLER_79_564 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2837 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xshift_reg_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2731 shift_reg_q\[15\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[11\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[11\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xrebuffer19 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ net51 VPWR VGND sg13g2_buf_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.sb_q\[14\] net2949 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2354 net1131 net2453 net2251 VPWR VGND sg13g2_a22oi_1
XFILLER_63_943 VPWR VGND sg13g2_fill_1
XFILLER_62_420 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[66\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2485 i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nor3_1_A_Y net2451 net2783 i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_dfrbpq_1_Q_D
+ net2912 sg13g2_a221oi_1
XFILLER_35_656 VPWR VGND sg13g2_fill_2
XFILLER_50_604 VPWR VGND sg13g2_fill_1
XFILLER_23_807 VPWR VGND sg13g2_fill_2
XFILLER_15_380 VPWR VGND sg13g2_decap_8
XFILLER_16_892 VPWR VGND sg13g2_fill_2
XFILLER_22_339 VPWR VGND sg13g2_fill_1
XFILLER_30_383 VPWR VGND sg13g2_decap_8
XFILLER_31_895 VPWR VGND sg13g2_fill_2
Xrsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1263 net3066 rsp_data_q\[0\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VGND net2568 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[275\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xhold502 strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B VPWR
+ VGND net534 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[94\]
+ net2843 i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
Xhold513 i_snitch.wake_up_q\[2\] VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold524 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold535 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net567 sg13g2_dlygate4sd3_1
XFILLER_103_105 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q
+ net3248 VGND VPWR net1086 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
Xhold546 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net578 sg13g2_dlygate4sd3_1
Xhold579 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net611 sg13g2_dlygate4sd3_1
Xhold568 i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y VPWR VGND net600 sg13g2_dlygate4sd3_1
Xhold557 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\] VPWR
+ VGND net589 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_100_812 VPWR VGND sg13g2_decap_8
XFILLER_58_748 VPWR VGND sg13g2_fill_2
Xhold1213 i_snitch.gpr_waddr\[4\] VPWR VGND net1245 sg13g2_dlygate4sd3_1
Xhold1202 i_snitch.i_snitch_regfile.mem\[123\] VPWR VGND net1234 sg13g2_dlygate4sd3_1
Xhold1224 i_snitch.i_snitch_lsu.metadata_q\[1\] VPWR VGND net1256 sg13g2_dlygate4sd3_1
XFILLER_73_718 VPWR VGND sg13g2_decap_4
Xhold1235 i_snitch.i_snitch_regfile.mem\[509\] VPWR VGND net1267 sg13g2_dlygate4sd3_1
Xhold1246 i_snitch.i_snitch_regfile.mem\[187\] VPWR VGND net1278 sg13g2_dlygate4sd3_1
Xhold1257 i_snitch.i_snitch_regfile.mem\[131\] VPWR VGND net1289 sg13g2_dlygate4sd3_1
XFILLER_100_889 VPWR VGND sg13g2_decap_8
Xhold1268 rsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1300 sg13g2_dlygate4sd3_1
XFILLER_66_781 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_26_612 VPWR VGND sg13g2_fill_1
Xhold1279 i_snitch.i_snitch_regfile.mem\[323\] VPWR VGND net1311 sg13g2_dlygate4sd3_1
XFILLER_39_984 VPWR VGND sg13g2_fill_2
XFILLER_25_122 VPWR VGND sg13g2_decap_8
XFILLER_81_762 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1
+ i_req_arb.data_i\[44\]_sg13g2_a21o_1_B1_X VPWR VGND sg13g2_nand2_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_41_604 VPWR VGND sg13g2_fill_2
XFILLER_90_1022 VPWR VGND sg13g2_decap_8
XFILLER_13_328 VPWR VGND sg13g2_decap_4
XFILLER_15_67 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B_sg13g2_nor4_1_Y
+ net3076 net3080 net3081 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ VGND VPWR net3075 sg13g2_nor4_2
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
Xrsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_snitch.sb_q\[11\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.sb_d\[11\] i_snitch.sb_q\[11\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xoutput22 net22 uo_out[5] VPWR VGND sg13g2_buf_1
Xoutput9 net9 uio_out[0] VPWR VGND sg13g2_buf_1
Xoutput11 net11 uio_out[2] VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A
+ i_snitch.inst_addr_o\[12\] net2527 VPWR VGND sg13g2_nand2_1
XFILLER_1_755 VPWR VGND sg13g2_decap_8
XFILLER_89_895 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X net2301 net1119 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[3\] VPWR VGND sg13g2_a21o_1
XFILLER_49_759 VPWR VGND sg13g2_fill_2
Xdata_pdata\[2\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C net3149 data_pdata\[10\]_sg13g2_nor2b_1_A_Y
+ data_pdata\[2\]_sg13g2_nor2_1_B_Y data_pdata\[2\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_102_182 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y
+ net3176 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_91_515 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_91_548 VPWR VGND sg13g2_fill_2
XFILLER_17_645 VPWR VGND sg13g2_fill_2
XFILLER_29_483 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[295\] clknet_leaf_117_clk sg13g2_dfrbpq_1
XFILLER_32_659 VPWR VGND sg13g2_fill_2
XFILLER_8_321 VPWR VGND sg13g2_fill_2
XFILLER_12_372 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2445 net2885 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
XFILLER_40_670 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[345\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2580 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_8_398 VPWR VGND sg13g2_fill_1
XFILLER_101_609 VPWR VGND sg13g2_decap_8
XFILLER_97_70 VPWR VGND sg13g2_decap_8
XFILLER_100_119 VPWR VGND sg13g2_decap_8
XFILLER_95_854 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[219\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net984 net2439 net2252 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_nand2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2827
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0 net3117 i_snitch.i_snitch_regfile.mem\[133\]
+ i_snitch.i_snitch_regfile.mem\[165\] i_snitch.i_snitch_regfile.mem\[197\] i_snitch.i_snitch_regfile.mem\[229\]
+ net3099 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_67_589 VPWR VGND sg13g2_fill_1
XFILLER_55_729 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ net2480 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ net2498 VPWR VGND sg13g2_a22oi_1
XFILLER_39_269 VPWR VGND sg13g2_decap_8
XFILLER_82_559 VPWR VGND sg13g2_decap_8
XFILLER_47_291 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[114\] clknet_leaf_88_clk sg13g2_dfrbpq_1
XFILLER_62_261 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q_D VGND net2329 net2257
+ sg13g2_o21ai_1
XFILLER_23_659 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2639 i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_50_478 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_11_1012 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[13\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net477 shift_reg_q\[13\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
XFILLER_105_959 VPWR VGND sg13g2_decap_8
Xhold398 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\] VPWR
+ VGND net430 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2419 sg13g2_a21oi_1
Xhold1010 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]
+ VPWR VGND net1042 sg13g2_dlygate4sd3_1
Xhold1021 i_snitch.i_snitch_regfile.mem\[39\] VPWR VGND net1053 sg13g2_dlygate4sd3_1
Xhold1032 i_snitch.i_snitch_regfile.mem\[231\] VPWR VGND net1064 sg13g2_dlygate4sd3_1
XFILLER_100_675 VPWR VGND sg13g2_fill_2
XFILLER_93_28 VPWR VGND sg13g2_decap_8
Xhold1076 rsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1108
+ sg13g2_dlygate4sd3_1
Xhold1054 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1086 sg13g2_dlygate4sd3_1
Xhold1043 i_snitch.inst_addr_o\[27\] VPWR VGND net1075 sg13g2_dlygate4sd3_1
Xhold1065 i_snitch.i_snitch_regfile.mem\[139\] VPWR VGND net1097 sg13g2_dlygate4sd3_1
XFILLER_39_781 VPWR VGND sg13g2_fill_2
Xhold1087 i_req_arb.data_i\[38\] VPWR VGND net1119 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2254 net2387 net1262 VPWR VGND sg13g2_a22oi_1
XFILLER_26_431 VPWR VGND sg13g2_decap_4
Xhold1098 i_snitch.i_snitch_regfile.mem\[398\] VPWR VGND net1130 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3170 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ state sg13g2_a21oi_1
XFILLER_42_957 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2720 i_snitch.inst_addr_o\[26\] sg13g2_a21oi_2
XFILLER_42_968 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
Xrsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1388 net3067 net1343 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1
+ net2555 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_101_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[239\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2333 net1128 net2677 net2877 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2641 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B net3163 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X VPWR VGND sg13g2_and2_1
XFILLER_104_970 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ net2523 VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.inst_addr_o\[27\] i_snitch.inst_addr_o\[28\] sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[134\] clknet_leaf_78_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_o21ai_1_A1 net2938 VPWR i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[301\] net2812 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3092 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_97_1006 VPWR VGND sg13g2_decap_8
XFILLER_92_813 VPWR VGND sg13g2_decap_4
XFILLER_76_386 VPWR VGND sg13g2_fill_1
XFILLER_76_375 VPWR VGND sg13g2_decap_4
XFILLER_36_206 VPWR VGND sg13g2_decap_4
XFILLER_92_857 VPWR VGND sg13g2_decap_8
XFILLER_91_323 VPWR VGND sg13g2_fill_2
XFILLER_76_397 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A_Y net2998 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net3027 sg13g2_a21oi_1
XFILLER_17_442 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y
+ VPWR VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X
+ sg13g2_nand4_1
XFILLER_72_570 VPWR VGND sg13g2_fill_1
XFILLER_44_261 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2711 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0 net3126 i_snitch.i_snitch_regfile.mem\[414\]
+ i_snitch.i_snitch_regfile.mem\[446\] i_snitch.i_snitch_regfile.mem\[478\] i_snitch.i_snitch_regfile.mem\[510\]
+ net3106 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_20_607 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[1\]_sg13g2_a22oi_1_A1 uio_out_sg13g2_inv_1_Y_2_A shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1_X
+ cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 shift_reg_q\[1\] VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[20\]_sg13g2_a21oi_1_A2 VGND VPWR net3160 data_pdata\[20\] data_pdata\[20\]_sg13g2_a21oi_1_A2_Y
+ net3153 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2386
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2704 i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_8_184 VPWR VGND sg13g2_decap_8
XFILLER_59_309 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2866
+ net2662 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[418\]_sg13g2_nor3_1_A net1339 net2865 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_67_320 VPWR VGND sg13g2_fill_1
XFILLER_55_504 VPWR VGND sg13g2_fill_2
XFILLER_103_49 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_83_879 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y VPWR
+ VGND sg13g2_nand2_2
XFILLER_23_401 VPWR VGND sg13g2_fill_2
XFILLER_24_935 VPWR VGND sg13g2_decap_4
XFILLER_11_607 VPWR VGND sg13g2_decap_8
XFILLER_23_467 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[154\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_o21ai_1_A1 net3107 VPWR i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[321\] net3128 sg13g2_o21ai_1
XFILLER_88_17 VPWR VGND sg13g2_decap_4
Xfanout3009 net3010 net3009 VPWR VGND sg13g2_buf_8
Xfanout2308 net2309 net2308 VPWR VGND sg13g2_buf_8
XFILLER_105_756 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2578 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xfanout2319 net2320 net2319 VPWR VGND sg13g2_buf_8
XFILLER_104_266 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B net3163 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[331\] VGND sg13g2_inv_1
XFILLER_101_973 VPWR VGND sg13g2_decap_8
XFILLER_74_835 VPWR VGND sg13g2_fill_1
XFILLER_18_228 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[18\] net854 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_14_445 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[103\]
+ net2998 i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_41_220 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2328
+ sg13g2_o21ai_1
XFILLER_6_611 VPWR VGND sg13g2_decap_4
XFILLER_6_644 VPWR VGND sg13g2_fill_1
XFILLER_6_699 VPWR VGND sg13g2_decap_8
Xfanout2820 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y
+ net2820 VPWR VGND sg13g2_buf_8
XFILLER_96_426 VPWR VGND sg13g2_fill_2
Xfanout2853 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B_X
+ net2853 VPWR VGND sg13g2_buf_8
XFILLER_78_83 VPWR VGND sg13g2_fill_1
Xdata_pdata\[16\]_sg13g2_nor2b_1_B_N net3159 data_pdata\[16\] data_pdata\[16\]_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_2_894 VPWR VGND sg13g2_decap_8
Xfanout2831 net2832 net2831 VPWR VGND sg13g2_buf_8
Xfanout2842 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y
+ net2842 VPWR VGND sg13g2_buf_8
Xfanout2864 net2865 net2864 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_2
Xfanout2897 data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2897 VPWR
+ VGND sg13g2_buf_8
Xfanout2886 net2887 net2886 VPWR VGND sg13g2_buf_8
Xfanout2875 net2877 net2875 VPWR VGND sg13g2_buf_8
XFILLER_76_161 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2325 net912 net2647 net2893 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C
+ net2640 i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_94_60 VPWR VGND sg13g2_fill_2
XFILLER_80_816 VPWR VGND sg13g2_decap_8
XFILLER_52_507 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR
+ VGND net2833 net2639 i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1_Y net2955
+ i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ sg13g2_a221oi_1
XFILLER_92_698 VPWR VGND sg13g2_fill_1
XFILLER_45_570 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[174\] clknet_leaf_88_clk sg13g2_dfrbpq_1
XFILLER_17_294 VPWR VGND sg13g2_fill_1
XFILLER_21_905 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1349 net2491 net1383 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3040
+ net2654 VPWR VGND sg13g2_nand2_1
Xdata_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2714 data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y
+ data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y net3070 sg13g2_a21oi_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_and3_1
XFILLER_101_203 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_and2_1_X
+ net116 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B
+ VPWR VGND sg13g2_and2_1
XFILLER_88_938 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[309\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_102_748 VPWR VGND sg13g2_decap_4
XFILLER_99_297 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_nor3_1
XFILLER_4_91 VPWR VGND sg13g2_decap_8
XFILLER_96_971 VPWR VGND sg13g2_decap_8
XFILLER_68_673 VPWR VGND sg13g2_decap_8
XFILLER_83_643 VPWR VGND sg13g2_decap_8
XFILLER_55_312 VPWR VGND sg13g2_decap_8
XFILLER_83_654 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2375 net881 net2651 net2743 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[116\]
+ net2806 i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_64_890 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2816 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2539 sg13g2_a21oi_1
XFILLER_23_264 VPWR VGND sg13g2_decap_8
XFILLER_51_584 VPWR VGND sg13g2_fill_1
XFILLER_8_909 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2702 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
XFILLER_99_49 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1369 net3066 net7 VPWR VGND sg13g2_a22oi_1
Xuo_out_sg13g2_buf_1_X_1 net3064 net18 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[299\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2680 net2780 net2318 net1351 VPWR VGND sg13g2_a22oi_1
XFILLER_2_102 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2919
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[361\]_sg13g2_o21ai_1_A1 net2969 VPWR i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[361\] net2802 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[194\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_93_407 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[500\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_19_515 VPWR VGND sg13g2_decap_8
XFILLER_87_993 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_46_334 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2862
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_104_70 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_0_49 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3084 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2849 net3075 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2751 sg13g2_a221oi_1
XFILLER_73_164 VPWR VGND sg13g2_fill_1
XFILLER_64_41 VPWR VGND sg13g2_fill_2
XFILLER_15_710 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[42\] clknet_leaf_94_clk sg13g2_dfrbpq_1
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_70_893 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[329\] clknet_leaf_50_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[118\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net982 net2651 net2871 VPWR VGND sg13g2_a22oi_1
Xhold909 data_pdata\[27\] VPWR VGND net941 sg13g2_dlygate4sd3_1
XFILLER_6_430 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2581 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net2578 sg13g2_a21oi_1
XFILLER_7_997 VPWR VGND sg13g2_decap_8
XFILLER_89_93 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2768
+ net2693 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ sg13g2_o21ai_1
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2459 net2283 net2369 net1241 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_o21ai_1_A1 net3013 VPWR i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[38\] net2990 sg13g2_o21ai_1
XFILLER_69_437 VPWR VGND sg13g2_fill_1
Xfanout2672 data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2672 VPWR VGND sg13g2_buf_8
Xfanout2661 net2662 net2661 VPWR VGND sg13g2_buf_8
XFILLER_2_691 VPWR VGND sg13g2_decap_8
Xfanout2650 data_pdata\[30\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2650 VPWR
+ VGND sg13g2_buf_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ net89 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X net2312 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1 VPWR VGND sg13g2_and2_1
Xfanout2683 i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N_Y
+ net2683 VPWR VGND sg13g2_buf_2
Xfanout2694 data_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2694 VPWR VGND sg13g2_buf_8
XFILLER_93_930 VPWR VGND sg13g2_decap_8
XFILLER_65_621 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
Xshift_reg_q\[17\]_sg13g2_a22oi_1_A1 shift_reg_q\[17\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_1_X
+ net3053 net3043 shift_reg_q\[17\] VPWR VGND sg13g2_a22oi_1
XFILLER_37_323 VPWR VGND sg13g2_fill_1
XFILLER_38_857 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q
+ net3203 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2878
+ net2674 VPWR VGND sg13g2_nand2_1
XFILLER_80_635 VPWR VGND sg13g2_fill_2
XFILLER_64_186 VPWR VGND sg13g2_fill_2
XFILLER_100_28 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[491\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[491\]
+ net3135 i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_a21oi_1_A1_Y net2945 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2833
+ VPWR i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2738
+ net2657 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[381\]_sg13g2_o21ai_1_A1 net2970 VPWR i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[381\] net2804 sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A_sg13g2_and3_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A
+ net2924 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_and3_1
Xclkload60 VPWR clkload60/Y clknet_leaf_81_clk VGND sg13g2_inv_1
XFILLER_47_1000 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A_Y net2845 i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_88_713 VPWR VGND sg13g2_decap_8
XFILLER_0_639 VPWR VGND sg13g2_decap_8
XFILLER_87_256 VPWR VGND sg13g2_fill_2
XFILLER_75_418 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[62\] clknet_leaf_94_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_A1
+ net2303 i_snitch.pc_d\[26\] i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2 i_snitch.inst_addr_o\[16\] i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_68_481 VPWR VGND sg13g2_fill_1
XFILLER_44_805 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ net2684 net2746 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_84_996 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[349\] clknet_leaf_95_clk sg13g2_dfrbpq_1
XFILLER_71_646 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[310\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[310\]
+ net3020 i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_a21oi_1_A1_Y net2990 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net852 net2446 net2282 VPWR VGND sg13g2_a22oi_1
XFILLER_24_573 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2499 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_24_584 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_o21ai_1_A1 net3004 VPWR i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[58\] net2977 sg13g2_o21ai_1
XFILLER_11_278 VPWR VGND sg13g2_fill_1
XFILLER_50_76 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ sg13g2_nand4_1
XFILLER_4_934 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2452
+ net2514 net2902 net2784 VPWR VGND sg13g2_a22oi_1
XFILLER_3_433 VPWR VGND sg13g2_decap_4
XFILLER_3_422 VPWR VGND sg13g2_fill_1
XFILLER_105_350 VPWR VGND sg13g2_decap_8
XFILLER_79_702 VPWR VGND sg13g2_fill_2
XFILLER_67_908 VPWR VGND sg13g2_decap_8
XFILLER_3_499 VPWR VGND sg13g2_fill_2
XFILLER_94_727 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.inst_addr_o\[17\]
+ net2528 VPWR VGND sg13g2_xnor2_1
XFILLER_66_418 VPWR VGND sg13g2_fill_2
XFILLER_75_941 VPWR VGND sg13g2_fill_1
XFILLER_19_356 VPWR VGND sg13g2_decap_8
Xdata_pdata\[3\]_sg13g2_dfrbpq_1_Q net3202 VGND VPWR net689 data_pdata\[3\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_B_N
+ VGND i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ sg13g2_o21ai_1
XFILLER_75_996 VPWR VGND sg13g2_fill_1
XFILLER_74_462 VPWR VGND sg13g2_fill_2
XFILLER_90_966 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C
+ net2421 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y VPWR VGND
+ sg13g2_nand2_1
XFILLER_62_646 VPWR VGND sg13g2_fill_2
Xdata_pdata\[5\]_sg13g2_mux2_1_A1 rsp_data_q\[5\] net676 net3048 data_pdata\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_34_326 VPWR VGND sg13g2_fill_2
XFILLER_61_145 VPWR VGND sg13g2_fill_1
XFILLER_43_860 VPWR VGND sg13g2_fill_2
Xrsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1223 net3064 rsp_data_q\[7\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[82\] clknet_leaf_87_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND net2783 sg13g2_nand2b_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
Xhold706 i_snitch.i_snitch_regfile.mem\[137\] VPWR VGND net738 sg13g2_dlygate4sd3_1
Xhold728 i_snitch.i_snitch_regfile.mem\[392\] VPWR VGND net760 sg13g2_dlygate4sd3_1
XFILLER_6_260 VPWR VGND sg13g2_fill_1
Xhold717 data_pdata\[18\] VPWR VGND net749 sg13g2_dlygate4sd3_1
Xhold739 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net771 sg13g2_dlygate4sd3_1
XFILLER_97_543 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_nand3b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y
+ VPWR VGND sg13g2_a22oi_1
Xfanout3181 net3181 net3182 VPWR VGND sg13g2_buf_16
Xfanout3170 net3171 net3170 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[369\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xfanout3192 net3193 net3192 VPWR VGND sg13g2_buf_8
Xfanout2480 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y
+ net2480 VPWR VGND sg13g2_buf_2
XFILLER_84_226 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net971 net2446 net2244 VPWR VGND sg13g2_a22oi_1
Xfanout2491 net2492 net2491 VPWR VGND sg13g2_buf_8
XFILLER_81_900 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_80_410 VPWR VGND sg13g2_decap_8
XFILLER_77_1026 VPWR VGND sg13g2_fill_2
XFILLER_53_602 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y
+ net2565 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_nor3_1
XFILLER_25_348 VPWR VGND sg13g2_fill_1
XFILLER_81_977 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2 VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_A1
+ i_snitch.pc_d\[8\] i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_Y i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y
+ net2745 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_576 VPWR VGND sg13g2_fill_2
XFILLER_4_219 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[336\] VGND sg13g2_inv_1
XFILLER_106_147 VPWR VGND sg13g2_decap_8
XFILLER_105_7 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_mux2_1_A1
+ net471 net609 net2617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.inst_addr_o\[29\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[29\]
+ i_snitch.inst_addr_o\[29\] clknet_leaf_54_clk sg13g2_dfrbpq_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_nand2_1_A_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_A2 net2623 sg13g2_o21ai_1
XFILLER_96_28 VPWR VGND sg13g2_decap_8
XFILLER_0_414 VPWR VGND sg13g2_decap_8
XFILLER_0_425 VPWR VGND sg13g2_fill_2
XFILLER_1_937 VPWR VGND sg13g2_decap_8
XFILLER_103_865 VPWR VGND sg13g2_decap_8
XFILLER_102_364 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1_X
+ VPWR VGND sg13g2_nand2b_1
XFILLER_29_632 VPWR VGND sg13g2_fill_1
Xdata_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR net3149 data_pdata\[19\]_sg13g2_mux2_1_A0_X
+ data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y data_pdata\[3\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_X
+ net3091 net2929 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_16_315 VPWR VGND sg13g2_fill_1
XFILLER_17_816 VPWR VGND sg13g2_fill_2
XFILLER_17_827 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1
+ net2561 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ net2579 sg13g2_o21ai_1
XFILLER_71_410 VPWR VGND sg13g2_fill_1
XFILLER_16_359 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_117_clk clknet_5_4__leaf_clk clknet_leaf_117_clk VPWR VGND sg13g2_buf_8
XFILLER_8_503 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_inv_1_A
+ net931 i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_A2 VPWR VGND sg13g2_inv_4
XFILLER_8_558 VPWR VGND sg13g2_fill_1
XFILLER_8_547 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[389\] clknet_leaf_110_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[178\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2444 net2272 net2344 net1178 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2533 net2419 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2500 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ VGND net2572 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_3_252 VPWR VGND sg13g2_fill_2
XFILLER_6_1019 VPWR VGND sg13g2_decap_8
XFILLER_67_749 VPWR VGND sg13g2_fill_1
XFILLER_66_204 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_39_418 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2
+ VGND VPWR net2546 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
XFILLER_75_771 VPWR VGND sg13g2_fill_1
XFILLER_90_763 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 net2489 sg13g2_o21ai_1
XFILLER_37_1010 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2632 VPWR i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_50_638 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_108_clk clknet_5_18__leaf_clk clknet_leaf_108_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ net2510 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_o21ai_1_A1_Y net3090 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q net3289 VGND VPWR i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[208\] clknet_leaf_89_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1 VPWR VGND
+ net2933 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y net3089 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold514 shift_reg_q\[16\] VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold536 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\] VPWR
+ VGND net568 sg13g2_dlygate4sd3_1
Xhold503 shift_reg_q\[1\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold525 i_snitch.sb_q\[13\] VPWR VGND net557 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A_sg13g2_nor4_1_Y
+ net2608 net2593 net2561 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ VGND VPWR net2589 sg13g2_nor4_2
Xhold547 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\] VPWR
+ VGND net579 sg13g2_dlygate4sd3_1
Xhold558 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net590 sg13g2_dlygate4sd3_1
Xhold569 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\] VPWR
+ VGND net601 sg13g2_dlygate4sd3_1
XFILLER_106_49 VPWR VGND sg13g2_decap_8
XFILLER_98_885 VPWR VGND sg13g2_decap_8
XFILLER_97_395 VPWR VGND sg13g2_fill_1
Xhold1203 i_req_arb.data_i\[40\] VPWR VGND net1235 sg13g2_dlygate4sd3_1
Xhold1214 i_snitch.i_snitch_regfile.mem\[312\] VPWR VGND net1246 sg13g2_dlygate4sd3_1
XFILLER_57_204 VPWR VGND sg13g2_decap_8
Xhold1225 i_snitch.i_snitch_regfile.mem\[298\] VPWR VGND net1257 sg13g2_dlygate4sd3_1
XFILLER_100_868 VPWR VGND sg13g2_decap_8
Xhold1236 i_snitch.i_snitch_regfile.mem\[313\] VPWR VGND net1268 sg13g2_dlygate4sd3_1
Xhold1247 i_snitch.i_snitch_regfile.mem\[35\] VPWR VGND net1279 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold1258 i_snitch.i_snitch_regfile.mem\[164\] VPWR VGND net1290 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2502 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xhold1269 i_snitch.i_snitch_regfile.mem\[419\] VPWR VGND net1301 sg13g2_dlygate4sd3_1
XFILLER_81_741 VPWR VGND sg13g2_fill_2
XFILLER_65_270 VPWR VGND sg13g2_fill_1
XFILLER_54_966 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[370\]
+ net3129 i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_a21oi_1_A1_Y net2943 sg13g2_a21oi_1
XFILLER_90_1001 VPWR VGND sg13g2_decap_8
XFILLER_81_796 VPWR VGND sg13g2_fill_1
XFILLER_15_24 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[198\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2337 net1113 net2900 net2791 VPWR VGND sg13g2_a22oi_1
XFILLER_40_104 VPWR VGND sg13g2_fill_1
XFILLER_80_295 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1
+ VGND net2931 net70 sg13g2_o21ai_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1
+ net46 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[504\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2370 net868 net2665 net2857 VPWR VGND sg13g2_a22oi_1
XFILLER_22_874 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ VGND net1160 net2488 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1124 net2687 net2768 VPWR VGND sg13g2_a22oi_1
Xoutput23 net23 uo_out[6] VPWR VGND sg13g2_buf_1
Xoutput12 net12 uio_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_734 VPWR VGND sg13g2_decap_8
XFILLER_103_651 VPWR VGND sg13g2_decap_4
XFILLER_89_874 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_102_161 VPWR VGND sg13g2_decap_8
XFILLER_88_362 VPWR VGND sg13g2_decap_4
XFILLER_76_524 VPWR VGND sg13g2_fill_2
XFILLER_56_75 VPWR VGND sg13g2_decap_4
XFILLER_56_42 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[47\]
+ net2828 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y net2823 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[228\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_45_988 VPWR VGND sg13g2_decap_8
XFILLER_45_966 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_q\[5\]_sg13g2_dfrbpq_1_Q net3250 VGND VPWR i_snitch.sb_d\[5\] i_snitch.sb_q\[5\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_60_947 VPWR VGND sg13g2_fill_2
XFILLER_60_936 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
XFILLER_8_344 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1354 net3064 net5 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2445 net2885 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
XFILLER_95_800 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[71\] VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] net651 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2577 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_95_833 VPWR VGND sg13g2_decap_8
XFILLER_79_384 VPWR VGND sg13g2_fill_2
XFILLER_79_373 VPWR VGND sg13g2_fill_2
XFILLER_94_321 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C net2518
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2 VPWR VGND sg13g2_nand3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_nand2_1_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_nand2_1_A_Y
+ net430 net2621 VPWR VGND sg13g2_nand2_1
XFILLER_48_760 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[322\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[280\]_sg13g2_o21ai_1_A1 net2938 VPWR i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[280\] i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_51_925 VPWR VGND sg13g2_fill_1
XFILLER_23_616 VPWR VGND sg13g2_decap_8
XFILLER_35_498 VPWR VGND sg13g2_fill_2
XFILLER_94_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2321
+ sg13g2_o21ai_1
XFILLER_16_690 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X
+ net2853 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1
+ VPWR VGND sg13g2_or3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2420 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_105_938 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2
+ VGND net2747 net47 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[248\] clknet_leaf_57_clk sg13g2_dfrbpq_1
Xhold399 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net431 sg13g2_dlygate4sd3_1
Xhold1000 i_snitch.i_snitch_regfile.mem\[233\] VPWR VGND net1032 sg13g2_dlygate4sd3_1
Xhold1033 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]
+ VPWR VGND net1065 sg13g2_dlygate4sd3_1
Xhold1011 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1043 sg13g2_dlygate4sd3_1
XFILLER_58_568 VPWR VGND sg13g2_decap_4
Xhold1022 data_pdata\[30\] VPWR VGND net1054 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\] net623 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_86_888 VPWR VGND sg13g2_decap_8
Xhold1066 i_snitch.i_snitch_regfile.mem\[157\] VPWR VGND net1098 sg13g2_dlygate4sd3_1
Xhold1055 i_snitch.i_snitch_regfile.mem\[149\] VPWR VGND net1087 sg13g2_dlygate4sd3_1
Xhold1044 i_snitch.i_snitch_regfile.mem\[50\] VPWR VGND net1076 sg13g2_dlygate4sd3_1
XFILLER_27_900 VPWR VGND sg13g2_decap_8
XFILLER_27_911 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2550 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
Xhold1077 i_snitch.i_snitch_regfile.mem\[502\] VPWR VGND net1109 sg13g2_dlygate4sd3_1
XFILLER_45_229 VPWR VGND sg13g2_decap_8
Xhold1088 i_snitch.i_snitch_regfile.mem\[476\] VPWR VGND net1120 sg13g2_dlygate4sd3_1
Xstrb_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2730 strb_reg_q\[1\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D strb_reg_q\[0\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold1099 i_snitch.i_snitch_regfile.mem\[93\] VPWR VGND net1131 sg13g2_dlygate4sd3_1
XFILLER_27_988 VPWR VGND sg13g2_fill_2
XFILLER_53_273 VPWR VGND sg13g2_decap_4
XFILLER_14_627 VPWR VGND sg13g2_decap_8
XFILLER_26_67 VPWR VGND sg13g2_fill_1
XFILLER_41_413 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ VGND sg13g2_inv_1
XFILLER_5_303 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2757 net2304
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2517 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_5_336 VPWR VGND sg13g2_decap_4
XFILLER_5_325 VPWR VGND sg13g2_decap_8
XFILLER_89_682 VPWR VGND sg13g2_fill_2
XFILLER_89_671 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_103_481 VPWR VGND sg13g2_fill_1
XFILLER_49_535 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[86\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net769 net2652 net2787 VPWR VGND sg13g2_a22oi_1
XFILLER_92_836 VPWR VGND sg13g2_decap_8
XFILLER_83_62 VPWR VGND sg13g2_fill_2
XFILLER_45_763 VPWR VGND sg13g2_fill_1
XFILLER_18_966 VPWR VGND sg13g2_fill_2
XFILLER_83_73 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2413
+ sg13g2_o21ai_1
XFILLER_32_402 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
XFILLER_60_799 VPWR VGND sg13g2_fill_2
XFILLER_13_693 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q net3308 VGND VPWR i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[268\] clknet_leaf_70_clk sg13g2_dfrbpq_1
XFILLER_8_163 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR net1105 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A_Y net3002 sg13g2_o21ai_1
XFILLER_99_424 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2496 i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_5_870 VPWR VGND sg13g2_fill_1
XFILLER_102_919 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_and2_1_B
+ net2591 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_80_1022 VPWR VGND sg13g2_decap_8
XFILLER_83_814 VPWR VGND sg13g2_decap_8
XFILLER_103_28 VPWR VGND sg13g2_decap_8
XFILLER_83_858 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[20\]_sg13g2_dfrbpq_1_Q net3231 VGND VPWR rsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[20\] clknet_leaf_30_clk sg13g2_dfrbpq_2
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[1\]_sg13g2_dfrbpq_1_Q net3235 VGND
+ VPWR net1399 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[1\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_82_368 VPWR VGND sg13g2_fill_2
XFILLER_91_891 VPWR VGND sg13g2_decap_8
XFILLER_51_711 VPWR VGND sg13g2_fill_2
XFILLER_36_785 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ net2549 VPWR VGND sg13g2_nand2_2
XFILLER_51_744 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2 VGND VPWR i_snitch.inst_addr_o\[25\]
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 sg13g2_a21oi_1
XFILLER_50_254 VPWR VGND sg13g2_fill_2
XFILLER_10_107 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_30_clk clknet_5_9__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
XFILLER_3_829 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B_sg13g2_nand3_1_Y
+ net2923 net2926 net3033 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_2_306 VPWR VGND sg13g2_fill_2
XFILLER_104_245 VPWR VGND sg13g2_decap_8
XFILLER_78_608 VPWR VGND sg13g2_fill_1
Xfanout2309 net2310 net2309 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2970 i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B_Y sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[13\] net1104 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ net3074 net2753 VPWR VGND sg13g2_nand2_2
XFILLER_101_952 VPWR VGND sg13g2_decap_8
XFILLER_98_490 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2573 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ net2539 sg13g2_a21oi_1
Xclkbuf_leaf_97_clk clknet_5_17__leaf_clk clknet_leaf_97_clk VPWR VGND sg13g2_buf_8
Xrsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ net1264 VGND sg13g2_inv_1
XFILLER_74_814 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_18_207 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q net3255 VGND VPWR i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[288\] clknet_leaf_106_clk sg13g2_dfrbpq_1
XFILLER_57_1024 VPWR VGND sg13g2_decap_4
XFILLER_15_969 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2416 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q
+ net3189 VGND VPWR net446 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
XFILLER_14_468 VPWR VGND sg13g2_fill_2
XFILLER_30_917 VPWR VGND sg13g2_fill_1
XFILLER_41_265 VPWR VGND sg13g2_fill_1
XFILLER_42_766 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_21_clk clknet_5_14__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_10_630 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2_1_A
+ net117 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ VPWR VGND sg13g2_nor2_2
XFILLER_5_144 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1_sg13g2_nand3_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ net2548 net2569 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1
+ VPWR VGND sg13g2_nand3_1
Xfanout2821 net2823 net2821 VPWR VGND sg13g2_buf_8
Xfanout2810 net2813 net2810 VPWR VGND sg13g2_buf_8
Xfanout2854 net2856 net2854 VPWR VGND sg13g2_buf_8
XFILLER_2_873 VPWR VGND sg13g2_decap_8
Xfanout2832 net2833 net2832 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[290\] VGND sg13g2_inv_1
Xfanout2843 net2847 net2843 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_88_clk clknet_5_21__leaf_clk clknet_leaf_88_clk VPWR VGND sg13g2_buf_8
Xfanout2865 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B_Y
+ net2865 VPWR VGND sg13g2_buf_8
Xfanout2876 net2877 net2876 VPWR VGND sg13g2_buf_8
Xfanout2887 net2890 net2887 VPWR VGND sg13g2_buf_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
Xfanout2898 data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2898 VPWR
+ VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2462 net2738 i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
XFILLER_64_313 VPWR VGND sg13g2_decap_4
XFILLER_92_677 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[107\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X
+ net3072 i_snitch.sb_q\[8\] i_snitch.sb_q\[9\] i_snitch.sb_q\[10\] i_snitch.sb_q\[11\]
+ net3071 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_mux4_1
XFILLER_18_730 VPWR VGND sg13g2_fill_1
XFILLER_33_722 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nand2b_1
XFILLER_91_198 VPWR VGND sg13g2_decap_4
XFILLER_72_390 VPWR VGND sg13g2_fill_1
XFILLER_45_593 VPWR VGND sg13g2_fill_1
XFILLER_33_755 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2481 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_12_clk clknet_5_3__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
XFILLER_9_494 VPWR VGND sg13g2_fill_2
XFILLER_9_483 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0 net3129 i_snitch.i_snitch_regfile.mem\[144\]
+ i_snitch.i_snitch_regfile.mem\[176\] i_snitch.i_snitch_regfile.mem\[208\] i_snitch.i_snitch_regfile.mem\[240\]
+ net3108 i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[98\]
+ net2800 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VGND i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X
+ sg13g2_o21ai_1
XFILLER_57_0 VPWR VGND sg13g2_decap_8
XFILLER_99_232 VPWR VGND sg13g2_decap_8
XFILLER_88_917 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2340
+ sg13g2_o21ai_1
XFILLER_102_716 VPWR VGND sg13g2_decap_4
XFILLER_99_287 VPWR VGND sg13g2_fill_1
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_96_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_79_clk clknet_5_28__leaf_clk clknet_leaf_79_clk VPWR VGND sg13g2_buf_8
XFILLER_101_259 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2357
+ sg13g2_o21ai_1
XFILLER_83_622 VPWR VGND sg13g2_decap_8
XFILLER_56_858 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2270 net2387 net1371 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[21\]_sg13g2_dfrbpq_1_Q net3191 VGND VPWR net804 data_pdata\[21\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y
+ VGND VPWR net2600 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_67_195 VPWR VGND sg13g2_fill_1
XFILLER_83_699 VPWR VGND sg13g2_decap_8
XFILLER_82_165 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2413
+ sg13g2_o21ai_1
XFILLER_63_390 VPWR VGND sg13g2_decap_4
XFILLER_51_563 VPWR VGND sg13g2_decap_4
XFILLER_24_788 VPWR VGND sg13g2_fill_2
XFILLER_99_28 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2544 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2611 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_20_983 VPWR VGND sg13g2_fill_1
XFILLER_87_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_mux4_1_A0 net3118 i_snitch.i_snitch_regfile.mem\[263\]
+ i_snitch.i_snitch_regfile.mem\[295\] i_snitch.i_snitch_regfile.mem\[327\] i_snitch.i_snitch_regfile.mem\[359\]
+ net3099 i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xuo_out_sg13g2_buf_1_X_2 strb_out net19 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[127\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_105_587 VPWR VGND sg13g2_fill_2
XFILLER_2_169 VPWR VGND sg13g2_fill_1
XFILLER_87_972 VPWR VGND sg13g2_decap_8
XFILLER_59_696 VPWR VGND sg13g2_decap_8
XFILLER_58_173 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[83\]
+ i_snitch.i_snitch_regfile.mem\[115\] net3120 i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ net95 i_snitch.inst_addr_o\[1\] i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ net2719 sg13g2_a221oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2
+ net45 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A VPWR
+ VGND sg13g2_a21o_2
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_19_549 VPWR VGND sg13g2_fill_1
XFILLER_62_839 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[26\]_sg13g2_dfrbpq_1_Q net3203 VGND VPWR net551 shift_reg_q\[26\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_64_86 VPWR VGND sg13g2_fill_2
XFILLER_15_755 VPWR VGND sg13g2_decap_4
XFILLER_27_593 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A
+ sg13g2_or2_1
XFILLER_70_872 VPWR VGND sg13g2_fill_2
XFILLER_15_799 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 VPWR VGND sg13g2_nand3_1
XFILLER_7_976 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ net2611 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[423\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2463 net2284 net2384 net1356 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ net2555 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2641 i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
Xfanout3330 rst_n net3330 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[327\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B
+ sg13g2_nor4_2
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_9_1006 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[354\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[354\] net3117 VPWR VGND sg13g2_nand2_1
XFILLER_97_758 VPWR VGND sg13g2_fill_1
Xfanout2651 net2652 net2651 VPWR VGND sg13g2_buf_8
XFILLER_2_670 VPWR VGND sg13g2_decap_8
Xfanout2662 data_pdata\[25\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2662 VPWR
+ VGND sg13g2_buf_8
Xfanout2640 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ net2640 VPWR VGND sg13g2_buf_8
Xfanout2684 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y
+ net2684 VPWR VGND sg13g2_buf_8
Xfanout2695 net2698 net2695 VPWR VGND sg13g2_buf_8
Xfanout2673 net2674 net2673 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_1_clk clknet_5_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_29_4 VPWR VGND sg13g2_decap_4
XFILLER_78_994 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2898 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VGND net2749 i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[86\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_nand2b_1_A_N_Y
+ net3029 i_snitch.i_snitch_regfile.mem\[86\] VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y
+ sg13g2_o21ai_1
XFILLER_93_986 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net2296 net1299 net2494 net1310 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[10\]_sg13g2_mux2_1_A1 rsp_data_q\[10\] net824 net3048 data_pdata\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_33_552 VPWR VGND sg13g2_fill_2
XFILLER_61_894 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q net3190 VGND VPWR i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[147\] clknet_leaf_122_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[314\] net2810 sg13g2_o21ai_1
Xrsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ net1224 VGND sg13g2_inv_1
XFILLER_106_329 VPWR VGND sg13g2_decap_8
Xclkload61 VPWR clkload61/Y clknet_leaf_61_clk VGND sg13g2_inv_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2773 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_2
Xclkload50 clknet_leaf_106_clk clkload50/X VPWR VGND sg13g2_buf_8
XFILLER_0_618 VPWR VGND sg13g2_decap_8
XFILLER_102_546 VPWR VGND sg13g2_decap_8
XFILLER_84_975 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2876
+ net2649 VPWR VGND sg13g2_nand2_1
XFILLER_18_46 VPWR VGND sg13g2_decap_4
XFILLER_93_1021 VPWR VGND sg13g2_decap_8
XFILLER_24_530 VPWR VGND sg13g2_decap_4
XFILLER_51_360 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[443\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2463 net2252 net2384 net1285 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ net47 sg13g2_or2_1
Xclkload0 clknet_5_7__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2470 VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2657 VPWR VGND sg13g2_nand2_1
XFILLER_106_885 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_3_467 VPWR VGND sg13g2_fill_2
XFILLER_79_758 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[444\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[444\]
+ net3012 i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_a21oi_1_A1_Y net2985 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2575 VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VGND i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2581 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ net2578 sg13g2_a21oi_1
XFILLER_62_603 VPWR VGND sg13g2_fill_1
XFILLER_47_677 VPWR VGND sg13g2_fill_2
XFILLER_46_176 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[167\] clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_90_945 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2772
+ net2669 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y net2840 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_61_168 VPWR VGND sg13g2_decap_4
XFILLER_98_7 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_decap_8
XFILLER_30_522 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1
+ net2307 i_snitch.pc_d\[30\] i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1 net2528 i_snitch.inst_addr_o\[18\] i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X VPWR VGND sg13g2_a21o_1
Xhold707 i_snitch.i_snitch_regfile.mem\[201\] VPWR VGND net739 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2654 VPWR VGND sg13g2_nand2_1
Xhold718 data_pdata\[18\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net750 sg13g2_dlygate4sd3_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C
+ VPWR VGND sg13g2_and4_1
Xhold729 i_snitch.i_snitch_regfile.mem\[255\] VPWR VGND net761 sg13g2_dlygate4sd3_1
XFILLER_97_511 VPWR VGND sg13g2_decap_8
Xfanout3182 net3182 net3183 VPWR VGND sg13g2_buf_16
Xfanout3171 net3172 net3171 VPWR VGND sg13g2_buf_8
Xfanout3160 net3161 net3160 VPWR VGND sg13g2_buf_2
XFILLER_3_990 VPWR VGND sg13g2_decap_8
XFILLER_85_706 VPWR VGND sg13g2_fill_2
Xfanout2481 net2483 net2481 VPWR VGND sg13g2_buf_8
Xfanout3193 net3194 net3193 VPWR VGND sg13g2_buf_8
Xfanout2470 net2471 net2470 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xfanout2492 net2493 net2492 VPWR VGND sg13g2_buf_8
XFILLER_38_611 VPWR VGND sg13g2_fill_1
XFILLER_84_249 VPWR VGND sg13g2_decap_8
XFILLER_65_430 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[463\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net744 net2677 net2741 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2573 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y
+ sg13g2_a21oi_1
XFILLER_93_761 VPWR VGND sg13g2_fill_1
XFILLER_77_1005 VPWR VGND sg13g2_decap_8
XFILLER_65_452 VPWR VGND sg13g2_fill_2
XFILLER_53_614 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y net3005 sg13g2_o21ai_1
XFILLER_92_293 VPWR VGND sg13g2_fill_1
XFILLER_81_956 VPWR VGND sg13g2_decap_8
XFILLER_65_485 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3172 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ state sg13g2_a21oi_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ net2593 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_33_371 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_126 VPWR VGND sg13g2_decap_8
Xtarget_sel_q_sg13g2_nand2b_1_A_N target_sel_q_sg13g2_nand2b_1_A_N_Y net914 VPWR VGND
+ target_sel_q sg13g2_nand2b_2
XFILLER_1_916 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0 net3001 i_snitch.i_snitch_regfile.mem\[389\]
+ i_snitch.i_snitch_regfile.mem\[421\] i_snitch.i_snitch_regfile.mem\[453\] i_snitch.i_snitch_regfile.mem\[485\]
+ net2974 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_103_844 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q net3192 VGND VPWR i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[187\] clknet_leaf_119_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[354\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[354\] net2801 sg13g2_o21ai_1
XFILLER_102_343 VPWR VGND sg13g2_decap_8
XFILLER_69_791 VPWR VGND sg13g2_fill_1
XFILLER_48_419 VPWR VGND sg13g2_decap_8
XFILLER_21_1015 VPWR VGND sg13g2_decap_8
XFILLER_83_260 VPWR VGND sg13g2_fill_1
XFILLER_83_282 VPWR VGND sg13g2_fill_1
XFILLER_43_102 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[35\] clknet_leaf_104_clk sg13g2_dfrbpq_1
XFILLER_71_444 VPWR VGND sg13g2_decap_8
XFILLER_25_861 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2712 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
Xdata_pdata\[17\]_sg13g2_mux2_1_A1 rsp_data_q\[17\] net729 net3052 data_pdata\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_40_820 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_o21ai_1_A2 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A
+ VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_o21ai_1_A2_Y VGND i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp
+ i_req_arb.gen_arbiter.req_d\[1\] sg13g2_o21ai_1
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
Xstrb_reg_q\[5\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net443 strb_reg_q\[5\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
XFILLER_6_49 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1271 net2495 net1230 VPWR VGND sg13g2_a22oi_1
XFILLER_4_743 VPWR VGND sg13g2_fill_1
XFILLER_79_500 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2738
+ net2661 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ sg13g2_a21oi_2
XFILLER_0_982 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q
+ net3199 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1_sg13g2_inv_1_Y
+ VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1
+ net2515 VGND sg13g2_inv_1
XFILLER_23_809 VPWR VGND sg13g2_fill_1
XFILLER_35_658 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[484\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[484\]
+ net3122 i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_a21oi_1_A1_Y net2946 sg13g2_a21oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N
+ VPWR VGND sg13g2_nand2b_1
XFILLER_16_894 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2735 shift_reg_q\[16\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[12\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[12\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_31_842 VPWR VGND sg13g2_fill_1
XFILLER_31_897 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[374\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[374\] net2808 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2782
+ net2898 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.data_o\[41\]_sg13g2_o21ai_1_Y i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.data_o\[41\] VGND net3164 i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xhold515 shift_reg_q\[16\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net547 sg13g2_dlygate4sd3_1
XFILLER_7_592 VPWR VGND sg13g2_decap_4
Xhold504 shift_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net536 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2687 net2779 net2317 net1231 VPWR VGND sg13g2_a22oi_1
Xhold526 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net558 sg13g2_dlygate4sd3_1
Xhold537 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\] VPWR
+ VGND net569 sg13g2_dlygate4sd3_1
Xhold548 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net580 sg13g2_dlygate4sd3_1
Xhold559 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\] VPWR
+ VGND net591 sg13g2_dlygate4sd3_1
Xdata_pdata\[21\]_sg13g2_mux2_1_A0 data_pdata\[21\] data_pdata\[29\] net3155 data_pdata\[21\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[55\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_106_28 VPWR VGND sg13g2_decap_8
XFILLER_98_864 VPWR VGND sg13g2_decap_8
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_97_363 VPWR VGND sg13g2_fill_1
Xhold1204 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\] VPWR
+ VGND net1236 sg13g2_dlygate4sd3_1
Xhold1215 i_snitch.i_snitch_regfile.mem\[132\] VPWR VGND net1247 sg13g2_dlygate4sd3_1
XFILLER_100_847 VPWR VGND sg13g2_decap_8
Xhold1237 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\] VPWR
+ VGND net1269 sg13g2_dlygate4sd3_1
Xhold1248 i_snitch.i_snitch_regfile.mem\[297\] VPWR VGND net1280 sg13g2_dlygate4sd3_1
Xhold1226 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] VPWR
+ VGND net1258 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
XFILLER_66_783 VPWR VGND sg13g2_fill_1
XFILLER_66_761 VPWR VGND sg13g2_decap_8
Xhold1259 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] VPWR
+ VGND net1291 sg13g2_dlygate4sd3_1
XFILLER_54_923 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_o21ai_1_A1 net2963 VPWR i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[509\] net2804 sg13g2_o21ai_1
XFILLER_38_452 VPWR VGND sg13g2_decap_4
XFILLER_39_986 VPWR VGND sg13g2_fill_1
XFILLER_65_260 VPWR VGND sg13g2_decap_4
XFILLER_25_102 VPWR VGND sg13g2_decap_4
XFILLER_14_809 VPWR VGND sg13g2_fill_2
XFILLER_25_157 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_fill_1
XFILLER_31_68 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xoutput24 net24 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput13 net13 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_713 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1
+ net1018 net642 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_89_853 VPWR VGND sg13g2_decap_8
XFILLER_0_223 VPWR VGND sg13g2_decap_8
XFILLER_102_140 VPWR VGND sg13g2_decap_8
XFILLER_0_278 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_76_547 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y sg13g2_o21ai_1
XFILLER_17_625 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C
+ net3147 net3142 VPWR VGND sg13g2_nand2b_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X
+ VPWR i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2958
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2970
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[75\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_nor3_1_A net1326 net2765 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
XFILLER_98_105 VPWR VGND sg13g2_decap_4
XFILLER_95_812 VPWR VGND sg13g2_fill_2
XFILLER_67_547 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]_sg13g2_nand2_1_B
+ i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_B1 net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[44\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_889 VPWR VGND sg13g2_decap_8
XFILLER_82_517 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A_sg13g2_nand2b_1_Y i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A
+ net2515 i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y VPWR VGND sg13g2_nand2b_1
XFILLER_54_219 VPWR VGND sg13g2_decap_4
XFILLER_36_945 VPWR VGND sg13g2_fill_2
XFILLER_90_572 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2816 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_22_138 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_105_917 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2479 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2530 VPWR VGND sg13g2_a22oi_1
XFILLER_104_427 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_633 VPWR VGND sg13g2_decap_8
XFILLER_86_867 VPWR VGND sg13g2_decap_8
Xhold1023 data_pdata\[30\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net1055 sg13g2_dlygate4sd3_1
Xhold1001 i_snitch.i_snitch_regfile.mem\[147\] VPWR VGND net1033 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[281\] VGND sg13g2_inv_1
Xhold1012 i_snitch.i_snitch_regfile.mem\[461\] VPWR VGND net1044 sg13g2_dlygate4sd3_1
XFILLER_85_355 VPWR VGND sg13g2_fill_1
Xhold1034 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1066 sg13g2_dlygate4sd3_1
Xhold1056 i_snitch.i_snitch_regfile.mem\[120\] VPWR VGND net1088 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[342\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2403 net743 net2652 net2796 VPWR VGND sg13g2_a22oi_1
Xhold1045 i_snitch.i_snitch_regfile.mem\[384\] VPWR VGND net1077 sg13g2_dlygate4sd3_1
Xhold1067 i_snitch.i_snitch_regfile.mem\[474\] VPWR VGND net1099 sg13g2_dlygate4sd3_1
XFILLER_100_688 VPWR VGND sg13g2_decap_4
XFILLER_85_388 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ net1348 VGND sg13g2_inv_1
Xhold1089 i_snitch.i_snitch_regfile.mem\[396\] VPWR VGND net1121 sg13g2_dlygate4sd3_1
Xhold1078 i_snitch.i_snitch_regfile.mem\[90\] VPWR VGND net1110 sg13g2_dlygate4sd3_1
XFILLER_39_783 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[95\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_26_46 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B
+ net38 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_53_263 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2551 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
XFILLER_42_959 VPWR VGND sg13g2_fill_1
XFILLER_10_845 VPWR VGND sg13g2_fill_2
XFILLER_10_878 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[1\]_sg13g2_dfrbpq_1_Q net3239 VGND VPWR rsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[1\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2386
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y
+ net2717 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B VPWR
+ VGND sg13g2_nor2_1
XFILLER_3_28 VPWR VGND sg13g2_decap_8
Xhold890 i_snitch.i_snitch_regfile.mem\[113\] VPWR VGND net922 sg13g2_dlygate4sd3_1
XFILLER_1_587 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2757 net2303
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2517 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_67_42 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_91_325 VPWR VGND sg13g2_fill_1
XFILLER_76_399 VPWR VGND sg13g2_fill_1
XFILLER_29_271 VPWR VGND sg13g2_fill_1
XFILLER_83_30 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_455 VPWR VGND sg13g2_fill_2
XFILLER_60_712 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR net617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_34_1014 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] net591 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_142 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[362\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net930 net2470 net2282 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X
+ VPWR VGND sg13g2_and4_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A
+ net3078 net2753 VPWR VGND sg13g2_nand2_1
XFILLER_80_1001 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2516 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A
+ net2427 sg13g2_a21oi_1
Xi_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[1\] clknet_leaf_11_clk sg13g2_dfrbpq_2
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VGND net2749 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ sg13g2_o21ai_1
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
XFILLER_95_664 VPWR VGND sg13g2_fill_2
XFILLER_55_506 VPWR VGND sg13g2_fill_1
XFILLER_94_163 VPWR VGND sg13g2_decap_4
XFILLER_82_336 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_91_870 VPWR VGND sg13g2_decap_8
XFILLER_63_561 VPWR VGND sg13g2_fill_1
XFILLER_35_263 VPWR VGND sg13g2_fill_2
XFILLER_35_274 VPWR VGND sg13g2_fill_2
XFILLER_90_380 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2476 i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2469 net2879 i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q_D net2908
+ sg13g2_a221oi_1
Xi_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B net3071
+ i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_12_15 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net1053 net2454 net2285 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_104_224 VPWR VGND sg13g2_decap_8
XFILLER_59_812 VPWR VGND sg13g2_decap_4
XFILLER_58_300 VPWR VGND sg13g2_decap_4
XFILLER_101_931 VPWR VGND sg13g2_decap_8
XFILLER_86_631 VPWR VGND sg13g2_decap_4
XFILLER_59_856 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_dfrbpq_1_Q
+ net3203 VGND VPWR net599 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_1
XFILLER_82_881 VPWR VGND sg13g2_decap_8
XFILLER_26_252 VPWR VGND sg13g2_decap_8
XFILLER_14_447 VPWR VGND sg13g2_fill_1
XFILLER_41_222 VPWR VGND sg13g2_fill_1
XFILLER_53_55 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2397 net1125 net2470 net2245 VPWR VGND sg13g2_a22oi_1
XFILLER_10_675 VPWR VGND sg13g2_decap_4
XFILLER_6_624 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[28\] net806 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2328
+ sg13g2_o21ai_1
XFILLER_10_697 VPWR VGND sg13g2_fill_1
XFILLER_5_123 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A
+ net3088 net3094 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2
+ VPWR VGND sg13g2_nor2_2
XFILLER_5_178 VPWR VGND sg13g2_decap_4
XFILLER_2_852 VPWR VGND sg13g2_decap_8
Xfanout2800 net2801 net2800 VPWR VGND sg13g2_buf_8
Xfanout2811 net2813 net2811 VPWR VGND sg13g2_buf_8
XFILLER_97_929 VPWR VGND sg13g2_decap_8
Xfanout2833 i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_B1 net2833 VPWR
+ VGND sg13g2_buf_8
Xfanout2844 net2847 net2844 VPWR VGND sg13g2_buf_8
Xfanout2855 net2856 net2855 VPWR VGND sg13g2_buf_8
Xfanout2822 net2823 net2822 VPWR VGND sg13g2_buf_8
Xfanout2866 net2867 net2866 VPWR VGND sg13g2_buf_8
Xfanout2888 net2889 net2888 VPWR VGND sg13g2_buf_8
Xfanout2877 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1_X
+ net2877 VPWR VGND sg13g2_buf_8
XFILLER_92_601 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_49_355 VPWR VGND sg13g2_fill_1
Xfanout2899 net2900 net2899 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_mux2_1_A0
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\] net579 net2624
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_64_358 VPWR VGND sg13g2_fill_1
XFILLER_64_347 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1
+ VGND net2603 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2377
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[412\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net1071 net2454 net2253 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_mux2_1_A0_X net3100 net2824 i_snitch.i_snitch_regfile.mem\[59\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_17_285 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1 VPWR VGND net3106 net2822
+ i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[62\]
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1_Y net2827 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[201\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2339 net739 net2686 net2790 VPWR VGND sg13g2_a22oi_1
XFILLER_60_542 VPWR VGND sg13g2_fill_1
XFILLER_20_406 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2462 net2739 i_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
XFILLER_20_439 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_9_462 VPWR VGND sg13g2_fill_1
XFILLER_13_491 VPWR VGND sg13g2_decap_8
XFILLER_101_238 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_83_601 VPWR VGND sg13g2_fill_1
XFILLER_68_664 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2415 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_95_461 VPWR VGND sg13g2_decap_4
XFILLER_28_517 VPWR VGND sg13g2_fill_1
XFILLER_28_539 VPWR VGND sg13g2_decap_8
XFILLER_71_807 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D
+ net2923 net2926 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y
+ sg13g2_nand4_1
Xshift_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2732 shift_reg_q\[4\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[0\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xshift_reg_q\[3\]_sg13g2_dfrbpq_1_Q net3188 VGND VPWR net522 shift_reg_q\[3\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_104_1012 VPWR VGND sg13g2_decap_8
XFILLER_20_962 VPWR VGND sg13g2_decap_4
Xi_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y net1367
+ net2488 i_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 VPWR VGND
+ sg13g2_nor2_1
XFILLER_87_1007 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\] net587 net2618
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xuo_out_sg13g2_buf_1_X_3 i_req_register.data_o\[5\] net20 VPWR VGND sg13g2_buf_1
Xdata_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2 data_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ net3070 net2714 data_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_2_137 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[432\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_101_761 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VGND net2709 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
XFILLER_87_951 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1 VPWR VGND i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2834 i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_nand2b_1_A_N_Y i_snitch.i_snitch_regfile.mem\[64\]
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y net2842 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net977 net2678 net2787 VPWR VGND sg13g2_a22oi_1
XFILLER_74_634 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[221\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net1016 net2440 net2250 VPWR VGND sg13g2_a22oi_1
XFILLER_100_282 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ net2545 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ net2699 VPWR VGND sg13g2_a22oi_1
XFILLER_64_43 VPWR VGND sg13g2_fill_1
XFILLER_70_840 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2920
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
XFILLER_70_851 VPWR VGND sg13g2_fill_1
XFILLER_64_98 VPWR VGND sg13g2_fill_2
XFILLER_42_553 VPWR VGND sg13g2_fill_1
XFILLER_9_49 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_inv_1_A_Y net3091 net2918 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2825
+ sg13g2_a221oi_1
XFILLER_11_984 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nor2b_1_B_N i_snitch.i_snitch_lsu.metadata_q\[9\] data_pvalid
+ data_pvalid_sg13g2_nor2b_1_B_N_Y VPWR VGND sg13g2_nor2b_2
XFILLER_6_421 VPWR VGND sg13g2_fill_1
XFILLER_6_487 VPWR VGND sg13g2_fill_1
Xfanout3320 net3325 net3320 VPWR VGND sg13g2_buf_1
Xfanout2630 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B_Y
+ net2630 VPWR VGND sg13g2_buf_8
Xfanout2641 net2642 net2641 VPWR VGND sg13g2_buf_8
Xfanout2652 data_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2652 VPWR
+ VGND sg13g2_buf_8
Xfanout2663 data_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2663 VPWR
+ VGND sg13g2_buf_8
Xfanout2696 net2698 net2696 VPWR VGND sg13g2_buf_8
XFILLER_78_973 VPWR VGND sg13g2_decap_8
Xfanout2685 net2686 net2685 VPWR VGND sg13g2_buf_8
Xfanout2674 data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2674 VPWR VGND sg13g2_buf_8
Xrsp_data_q\[13\]_sg13g2_dfrbpq_1_Q net3239 VGND VPWR rsp_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[13\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_77_461 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_A1
+ net1405 VPWR VGND sg13g2_inv_2
XFILLER_93_965 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_65_656 VPWR VGND sg13g2_fill_2
XFILLER_92_464 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xnor2_1_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xnor2_1
XFILLER_53_829 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_nor3_1_A net1341 net3039 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B
+ net2763 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_64_188 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[304\] VGND sg13g2_inv_1
XFILLER_33_531 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2870
+ net2693 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[452\] clknet_leaf_109_clk sg13g2_dfrbpq_1
XFILLER_106_308 VPWR VGND sg13g2_decap_8
Xclkload62 VPWR clkload62/Y clknet_leaf_62_clk VGND sg13g2_inv_1
Xclkload51 VPWR clkload51/Y clknet_leaf_73_clk VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[286\] VGND sg13g2_inv_1
Xclkload40 clkload40/Y clknet_leaf_94_clk VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[241\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2333 net979 net2664 net2877 VPWR VGND sg13g2_a22oi_1
XFILLER_102_514 VPWR VGND sg13g2_decap_4
XFILLER_69_962 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[320\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[320\] net2949 VPWR VGND sg13g2_nand2_1
XFILLER_69_995 VPWR VGND sg13g2_decap_8
XFILLER_95_280 VPWR VGND sg13g2_fill_1
XFILLER_84_954 VPWR VGND sg13g2_decap_8
XFILLER_83_442 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y VGND VPWR net2760 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2 net2305 sg13g2_a21oi_1
XFILLER_55_133 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[448\]_sg13g2_o21ai_1_A1 net2962 VPWR i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[448\] i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
XFILLER_44_807 VPWR VGND sg13g2_fill_1
XFILLER_43_317 VPWR VGND sg13g2_fill_2
XFILLER_93_1000 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR net759 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_37_892 VPWR VGND sg13g2_decap_4
XFILLER_52_862 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2641 i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_54_1028 VPWR VGND sg13g2_fill_1
Xclkload1 clknet_5_15__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2627 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ net2758 VPWR VGND sg13g2_a22oi_1
XFILLER_4_969 VPWR VGND sg13g2_decap_8
XFILLER_106_864 VPWR VGND sg13g2_decap_8
XFILLER_79_726 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y_sg13g2_nand3_1_B
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_C
+ VPWR VGND sg13g2_nand3_1
XFILLER_105_385 VPWR VGND sg13g2_decap_8
XFILLER_94_718 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3080 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2850 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2753 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ net2725 net74 sg13g2_a21oi_2
XFILLER_101_580 VPWR VGND sg13g2_fill_1
XFILLER_86_280 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1 VPWR VGND
+ net3091 net2929 i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ sg13g2_a221oi_1
XFILLER_19_347 VPWR VGND sg13g2_decap_4
XFILLER_90_924 VPWR VGND sg13g2_decap_8
XFILLER_35_829 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3105 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ net2850 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2754 sg13g2_a221oi_1
XFILLER_62_648 VPWR VGND sg13g2_fill_1
XFILLER_46_199 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[472\] clknet_leaf_59_clk sg13g2_dfrbpq_1
Xdata_pdata\[15\]_sg13g2_nand2b_1_B data_pdata\[15\]_sg13g2_nand2b_1_B_Y data_pdata\[15\]
+ net3160 VPWR VGND sg13g2_nand2b_1
XFILLER_30_501 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1
+ net1395 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2446
+ net2513 net2901 net2888 VPWR VGND sg13g2_a22oi_1
Xhold719 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\] VPWR
+ VGND net751 sg13g2_dlygate4sd3_1
Xhold708 i_snitch.i_snitch_regfile.mem\[140\] VPWR VGND net740 sg13g2_dlygate4sd3_1
XFILLER_7_774 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B net2767 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1
+ net2506 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_2
XFILLER_97_534 VPWR VGND sg13g2_decap_8
Xfanout3183 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q net3183
+ VPWR VGND sg13g2_buf_8
Xfanout3172 net3173 net3172 VPWR VGND sg13g2_buf_8
Xfanout3161 net3162 net3161 VPWR VGND sg13g2_buf_1
Xfanout3150 net3151 net3150 VPWR VGND sg13g2_buf_8
Xfanout3194 net3226 net3194 VPWR VGND sg13g2_buf_8
Xfanout2460 net2462 net2460 VPWR VGND sg13g2_buf_8
Xfanout2471 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2471 VPWR
+ VGND sg13g2_buf_8
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1_X
+ VPWR VGND sg13g2_and2_1
Xfanout2482 net2483 net2482 VPWR VGND sg13g2_buf_1
Xdata_pdata\[14\]_sg13g2_dfrbpq_1_Q net3203 VGND VPWR net1036 data_pdata\[14\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
Xfanout2493 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_o21ai_1_A2_Y net2493 VPWR VGND
+ sg13g2_buf_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y
+ net2592 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_66_954 VPWR VGND sg13g2_fill_1
XFILLER_38_634 VPWR VGND sg13g2_fill_1
XFILLER_65_464 VPWR VGND sg13g2_decap_8
XFILLER_26_829 VPWR VGND sg13g2_fill_2
XFILLER_37_144 VPWR VGND sg13g2_fill_2
XFILLER_37_166 VPWR VGND sg13g2_decap_4
XFILLER_81_935 VPWR VGND sg13g2_decap_8
XFILLER_77_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[155\]
+ i_snitch.i_snitch_regfile.mem\[187\] i_snitch.i_snitch_regfile.mem\[219\] i_snitch.i_snitch_regfile.mem\[251\]
+ net3098 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net2962 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2
+ net3093 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2751 sg13g2_a221oi_1
Xi_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net3154 net2486 i_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_80_489 VPWR VGND sg13g2_decap_8
XFILLER_61_681 VPWR VGND sg13g2_decap_8
XFILLER_33_361 VPWR VGND sg13g2_fill_1
XFILLER_61_692 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_105 VPWR VGND sg13g2_decap_8
XFILLER_101_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1
+ net3071 VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2827
+ sg13g2_a221oi_1
XFILLER_103_823 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2792
+ net2653 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nand2b_1_A_N_Y
+ net3026 i_snitch.i_snitch_regfile.mem\[66\] VPWR VGND sg13g2_nand2b_1
XFILLER_102_322 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[492\] clknet_leaf_69_clk sg13g2_dfrbpq_1
Xi_req_arb.data_i\[39\]_sg13g2_dfrbpq_1_Q net3261 VGND VPWR i_snitch.pc_d\[4\] i_req_arb.data_i\[39\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_60_1021 VPWR VGND sg13g2_decap_8
XFILLER_102_399 VPWR VGND sg13g2_fill_2
XFILLER_75_239 VPWR VGND sg13g2_decap_8
XFILLER_57_943 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_a22oi_1_B2_Y
+ net2323 net700 net2433 net2267 VPWR VGND sg13g2_a22oi_1
XFILLER_28_100 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[19\]_sg13g2_dfrbpq_1_Q net3197 VGND VPWR net499 shift_reg_q\[19\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
XFILLER_28_155 VPWR VGND sg13g2_fill_1
XFILLER_72_946 VPWR VGND sg13g2_fill_2
XFILLER_71_434 VPWR VGND sg13g2_fill_2
XFILLER_71_423 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 VGND
+ sg13g2_inv_1
XFILLER_24_350 VPWR VGND sg13g2_fill_1
XFILLER_101_84 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2959
+ i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2966
+ i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
Xshift_reg_q\[12\]_sg13g2_nor2_1_A net548 net2735 shift_reg_q\[12\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_8_549 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ net2580 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[94\]
+ i_snitch.i_snitch_regfile.mem\[126\] net3127 i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[416\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2384 net886 net2903 net2861 VPWR VGND sg13g2_a22oi_1
XFILLER_3_243 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2464 VPWR VGND sg13g2_nand2_1
XFILLER_106_683 VPWR VGND sg13g2_decap_8
XFILLER_79_523 VPWR VGND sg13g2_fill_1
XFILLER_79_512 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q net3310 VGND VPWR i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[311\] clknet_leaf_69_clk sg13g2_dfrbpq_1
XFILLER_3_276 VPWR VGND sg13g2_fill_2
XFILLER_105_182 VPWR VGND sg13g2_decap_8
XFILLER_0_961 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A
+ net2601 VPWR VGND sg13g2_nand2_1
XFILLER_66_228 VPWR VGND sg13g2_decap_4
XFILLER_75_762 VPWR VGND sg13g2_fill_1
XFILLER_63_902 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0 net3123 i_snitch.i_snitch_regfile.mem\[393\]
+ i_snitch.i_snitch_regfile.mem\[425\] i_snitch.i_snitch_regfile.mem\[457\] i_snitch.i_snitch_regfile.mem\[489\]
+ net3103 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_47_475 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2788
+ net2897 VPWR VGND sg13g2_nand2_1
XFILLER_19_188 VPWR VGND sg13g2_fill_2
XFILLER_62_434 VPWR VGND sg13g2_decap_8
XFILLER_16_851 VPWR VGND sg13g2_fill_2
XFILLER_62_478 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[307\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[307\] net2810 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2873
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_42_180 VPWR VGND sg13g2_decap_8
Xhold527 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\] VPWR
+ VGND net559 sg13g2_dlygate4sd3_1
Xhold516 shift_reg_q\[12\] VPWR VGND net548 sg13g2_dlygate4sd3_1
XFILLER_7_582 VPWR VGND sg13g2_decap_4
Xhold505 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] VPWR
+ VGND net537 sg13g2_dlygate4sd3_1
Xhold549 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\] VPWR
+ VGND net581 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_a21o_2
Xdata_pdata\[21\]_sg13g2_mux2_1_A1 rsp_data_q\[21\] net803 net3049 data_pdata\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xhold538 i_snitch.sb_q\[9\] VPWR VGND net570 sg13g2_dlygate4sd3_1
XFILLER_103_119 VPWR VGND sg13g2_decap_8
XFILLER_98_843 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B_sg13g2_and4_1_X
+ net3034 net2924 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B
+ VPWR VGND sg13g2_and4_1
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_32_0 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2489 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_o21ai_1
Xshift_reg_q\[7\]_sg13g2_a22oi_1_A1 shift_reg_q\[7\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_1_X
+ net3055 net3045 net492 VPWR VGND sg13g2_a22oi_1
XFILLER_100_826 VPWR VGND sg13g2_decap_8
XFILLER_85_504 VPWR VGND sg13g2_fill_2
Xhold1216 i_snitch.i_snitch_regfile.mem\[496\] VPWR VGND net1248 sg13g2_dlygate4sd3_1
Xhold1205 i_snitch.i_snitch_regfile.mem\[68\] VPWR VGND net1237 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]
+ net3179 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xrsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_57_228 VPWR VGND sg13g2_decap_8
Xhold1227 i_snitch.i_snitch_regfile.mem\[179\] VPWR VGND net1259 sg13g2_dlygate4sd3_1
Xhold1238 i_snitch.i_snitch_regfile.mem\[450\] VPWR VGND net1270 sg13g2_dlygate4sd3_1
Xfanout2290 net2291 net2290 VPWR VGND sg13g2_buf_8
Xhold1249 i_snitch.i_snitch_regfile.mem\[452\] VPWR VGND net1281 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[446\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net454 net2383 VPWR VGND sg13g2_nand2_1
XFILLER_53_401 VPWR VGND sg13g2_decap_4
XFILLER_53_434 VPWR VGND sg13g2_fill_2
XFILLER_25_136 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1
+ net2748 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[436\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net1034 net2671 net2863 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1345 net2492 net1265 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_21_331 VPWR VGND sg13g2_decap_8
XFILLER_21_342 VPWR VGND sg13g2_fill_1
XFILLER_22_876 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[25\]_sg13g2_nor2_1_A net515 net2728 shift_reg_q\[25\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[331\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_or2_1_X
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A
+ net3087 net3085 sg13g2_or2_1
XFILLER_31_36 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_a221oi_1_B1
+ VPWR VGND i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net1088 net2665 net2871 VPWR VGND sg13g2_a22oi_1
Xoutput14 net14 uio_out[5] VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_o21ai_1_A1 net3019 VPWR i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[40\] net2982 sg13g2_o21ai_1
XFILLER_0_202 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_1_769 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y net1392 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B
+ i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y net3009 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2657 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_102_196 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2660 VPWR VGND sg13g2_nand2_1
XFILLER_45_902 VPWR VGND sg13g2_fill_2
XFILLER_29_453 VPWR VGND sg13g2_fill_1
XFILLER_57_795 VPWR VGND sg13g2_fill_1
XFILLER_56_261 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_o21ai_1_A2
+ net3054 VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ VGND net3167 net471 sg13g2_o21ai_1
XFILLER_60_905 VPWR VGND sg13g2_decap_4
XFILLER_72_798 VPWR VGND sg13g2_fill_1
XFILLER_71_253 VPWR VGND sg13g2_fill_2
XFILLER_16_158 VPWR VGND sg13g2_fill_1
XFILLER_25_692 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_331 VPWR VGND sg13g2_fill_1
XFILLER_8_313 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2546 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2
+ net2957 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2962 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C_Y VPWR
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N_Y
+ sg13g2_nand4_1
XFILLER_99_629 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D
+ sg13g2_nor4_2
XFILLER_97_84 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xnor2_1
XFILLER_79_375 VPWR VGND sg13g2_fill_1
XFILLER_67_504 VPWR VGND sg13g2_fill_2
XFILLER_95_868 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[456\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net815 net2644 net2741 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2464
+ net2262 net2667 net2862 VPWR VGND sg13g2_a22oi_1
XFILLER_75_592 VPWR VGND sg13g2_fill_2
XFILLER_47_261 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[351\] clknet_leaf_70_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B_sg13g2_and3_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ i_req_arb.data_i\[43\] net3082 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X
+ VPWR VGND sg13g2_and3_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2708 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2553 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1_sg13g2_and3_1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1
+ net3033 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ VPWR VGND sg13g2_and3_1
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net740 net2692 net2888 VPWR VGND sg13g2_a22oi_1
XFILLER_16_692 VPWR VGND sg13g2_fill_1
XFILLER_22_128 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2782
+ net2662 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2501 net2422 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ sg13g2_a221oi_1
XFILLER_7_60 VPWR VGND sg13g2_decap_8
XFILLER_11_1026 VPWR VGND sg13g2_fill_2
XFILLER_104_406 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_B
+ net3147 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[347\] i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_645 VPWR VGND sg13g2_fill_2
XFILLER_86_846 VPWR VGND sg13g2_decap_8
XFILLER_85_334 VPWR VGND sg13g2_fill_1
XFILLER_85_323 VPWR VGND sg13g2_fill_2
Xhold1024 i_snitch.i_snitch_regfile.mem\[236\] VPWR VGND net1056 sg13g2_dlygate4sd3_1
Xhold1013 i_snitch.i_snitch_regfile.mem\[182\] VPWR VGND net1045 sg13g2_dlygate4sd3_1
Xhold1002 i_snitch.i_snitch_regfile.mem\[436\] VPWR VGND net1034 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B
+ net2958 i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xhold1057 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]
+ VPWR VGND net1089 sg13g2_dlygate4sd3_1
Xhold1046 i_snitch.i_snitch_regfile.mem\[183\] VPWR VGND net1078 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y net3133 sg13g2_o21ai_1
Xhold1035 i_snitch.i_snitch_regfile.mem\[284\] VPWR VGND net1067 sg13g2_dlygate4sd3_1
Xi_snitch.inst_addr_o\[11\]_sg13g2_dfrbpq_1_Q net3313 VGND VPWR i_snitch.pc_d\[11\]
+ i_snitch.inst_addr_o\[11\] clknet_leaf_55_clk sg13g2_dfrbpq_2
Xhold1079 i_snitch.i_snitch_regfile.mem\[404\] VPWR VGND net1111 sg13g2_dlygate4sd3_1
Xhold1068 i_snitch.i_snitch_regfile.mem\[406\] VPWR VGND net1100 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2574 VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VGND net2586 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xstrb_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2727 strb_reg_q\[2\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D strb_reg_q\[1\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_22_684 VPWR VGND sg13g2_fill_2
XFILLER_6_817 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net1120 net2461 net2247 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q
+ net3245 VGND VPWR net748 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
XFILLER_89_640 VPWR VGND sg13g2_decap_4
Xhold880 i_snitch.i_snitch_regfile.mem\[279\] VPWR VGND net912 sg13g2_dlygate4sd3_1
Xhold891 i_snitch.i_snitch_regfile.mem\[61\] VPWR VGND net923 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2478 i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2433 net2892 i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
XFILLER_104_984 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_77_824 VPWR VGND sg13g2_decap_8
Xdata_pdata\[28\]_sg13g2_mux2_1_A1 net1051 net1083 net3050 data_pdata\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_49_515 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[371\] clknet_leaf_115_clk sg13g2_dfrbpq_1
XFILLER_1_555 VPWR VGND sg13g2_fill_2
XFILLER_1_566 VPWR VGND sg13g2_decap_8
XFILLER_103_472 VPWR VGND sg13g2_fill_1
XFILLER_77_846 VPWR VGND sg13g2_fill_1
XFILLER_77_835 VPWR VGND sg13g2_fill_2
XFILLER_76_312 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q
+ net3230 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_67_65 VPWR VGND sg13g2_decap_8
XFILLER_49_537 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ VGND net2571 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_67_76 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[160\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2343 net910 net2903 net2773 VPWR VGND sg13g2_a22oi_1
XFILLER_18_902 VPWR VGND sg13g2_fill_2
XFILLER_32_404 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2761 net2309
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2519 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[367\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[367\] net2808 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2347
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[506\] clknet_leaf_116_clk sg13g2_dfrbpq_1
Xrsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_8_165 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N
+ net98 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2817 i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[48\] clknet_leaf_89_clk sg13g2_dfrbpq_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C
+ net99 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y
+ VPWR VGND i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N
+ sg13g2_nand4_1
Xi_snitch.inst_addr_o\[31\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[31\]
+ i_snitch.inst_addr_o\[31\] clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_4_382 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y net2717
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_51_713 VPWR VGND sg13g2_fill_1
XFILLER_35_242 VPWR VGND sg13g2_decap_8
Xcnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y
+ cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A VPWR VGND shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ sg13g2_nand2b_2
XFILLER_35_297 VPWR VGND sg13g2_fill_2
XFILLER_50_256 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[496\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2458 net2262 net2369 net1248 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_a21oi_1
XFILLER_10_109 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q net3211 VGND VPWR i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[391\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[180\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net866 net2671 net2775 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
XFILLER_104_203 VPWR VGND sg13g2_decap_8
XFILLER_2_308 VPWR VGND sg13g2_fill_1
XFILLER_101_910 VPWR VGND sg13g2_decap_8
XFILLER_99_993 VPWR VGND sg13g2_decap_8
XFILLER_59_846 VPWR VGND sg13g2_fill_1
XFILLER_86_665 VPWR VGND sg13g2_fill_1
XFILLER_59_879 VPWR VGND sg13g2_fill_1
XFILLER_101_987 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2
+ net2570 VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ VGND i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_96_1020 VPWR VGND sg13g2_decap_8
XFILLER_82_860 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[23\] net836 net2914 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[44\] VGND sg13g2_inv_1
XFILLER_54_562 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B
+ net120 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1 i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_Y
+ i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_Y i_req_arb.gen_arbiter.req_d\[1\] i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2
+ net763 VPWR VGND sg13g2_a22oi_1
XFILLER_53_45 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2430 net2253 net2316 net1162 VPWR VGND sg13g2_a22oi_1
XFILLER_14_415 VPWR VGND sg13g2_decap_8
XFILLER_14_426 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_41_256 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1_sg13g2_nand2_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[68\]_sg13g2_dfrbpq_1_Q net3224 VGND VPWR i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[68\] clknet_leaf_107_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[210\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_5_102 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2321
+ sg13g2_o21ai_1
Xuio_out_sg13g2_buf_1_X i_req_register.data_o\[42\] net13 VPWR VGND sg13g2_buf_1
XFILLER_97_908 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2515 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2427 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[277\] VGND sg13g2_inv_1
XFILLER_2_831 VPWR VGND sg13g2_decap_8
Xfanout2801 net2802 net2801 VPWR VGND sg13g2_buf_8
Xfanout2812 net2813 net2812 VPWR VGND sg13g2_buf_8
XFILLER_78_53 VPWR VGND sg13g2_fill_2
Xfanout2834 i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1_B1 net2834 VPWR
+ VGND sg13g2_buf_8
Xfanout2823 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a21oi_1_A1_B1 net2823 VPWR
+ VGND sg13g2_buf_8
Xfanout2845 net2846 net2845 VPWR VGND sg13g2_buf_8
XFILLER_104_781 VPWR VGND sg13g2_decap_8
XFILLER_77_621 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_fill_2
XFILLER_49_301 VPWR VGND sg13g2_fill_2
Xfanout2878 net2884 net2878 VPWR VGND sg13g2_buf_8
Xtarget_sel_q_sg13g2_dfrbpq_1_Q net3184 VGND VPWR net1027 target_sel_q clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
Xfanout2867 net2868 net2867 VPWR VGND sg13g2_buf_8
Xfanout2856 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y
+ net2856 VPWR VGND sg13g2_buf_8
XFILLER_103_280 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2334
+ sg13g2_o21ai_1
Xfanout2889 net2890 net2889 VPWR VGND sg13g2_buf_8
XFILLER_92_613 VPWR VGND sg13g2_fill_2
XFILLER_64_326 VPWR VGND sg13g2_fill_2
XFILLER_94_96 VPWR VGND sg13g2_fill_1
XFILLER_76_186 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3165 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ state sg13g2_a21oi_1
XFILLER_92_679 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2365
+ sg13g2_o21ai_1
XFILLER_17_264 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_72_381 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_32_212 VPWR VGND sg13g2_fill_1
XFILLER_32_223 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B_Y VPWR VGND
+ sg13g2_nor3_1
XFILLER_32_234 VPWR VGND sg13g2_fill_2
XFILLER_13_470 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X
+ net3033 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_and4_1
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y net2739 VPWR VGND sg13g2_nand2b_1
Xdata_pdata\[9\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net890 data_pdata\[9\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_9_496 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2481 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y
+ net2533 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ net2551 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_691 VPWR VGND sg13g2_fill_2
XFILLER_87_407 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_101_217 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]
+ net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_2
Xi_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 net2488 i_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_a22oi_1_B2_Y
+ net2404 net656 net2677 net2797 VPWR VGND sg13g2_a22oi_1
XFILLER_96_985 VPWR VGND sg13g2_decap_8
XFILLER_68_687 VPWR VGND sg13g2_decap_8
XFILLER_56_838 VPWR VGND sg13g2_decap_8
XFILLER_95_495 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[88\] clknet_leaf_59_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2701 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_83_679 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[230\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_23_223 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.inst_addr_o\[26\] net2524 VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1 net2527 VPWR VGND sg13g2_xnor2_1
XFILLER_23_48 VPWR VGND sg13g2_decap_8
XFILLER_105_512 VPWR VGND sg13g2_fill_1
XFILLER_105_501 VPWR VGND sg13g2_fill_1
Xuo_out_sg13g2_buf_1_X_4 i_req_register.data_o\[38\] net21 VPWR VGND sg13g2_buf_1
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_78_418 VPWR VGND sg13g2_decap_8
XFILLER_99_790 VPWR VGND sg13g2_decap_8
XFILLER_87_930 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2569 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
XFILLER_100_261 VPWR VGND sg13g2_decap_8
XFILLER_74_602 VPWR VGND sg13g2_decap_4
XFILLER_19_529 VPWR VGND sg13g2_fill_2
XFILLER_104_84 VPWR VGND sg13g2_decap_8
XFILLER_55_860 VPWR VGND sg13g2_fill_1
XFILLER_64_88 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2_B1_sg13g2_nor2b_1_Y
+ net3165 net666 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2_B1
+ VPWR VGND sg13g2_nor2b_1
XFILLER_54_392 VPWR VGND sg13g2_fill_2
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_30_738 VPWR VGND sg13g2_fill_1
XFILLER_80_76 VPWR VGND sg13g2_fill_1
XFILLER_10_440 VPWR VGND sg13g2_fill_2
Xfanout3321 net3325 net3321 VPWR VGND sg13g2_buf_8
Xfanout3310 net3311 net3310 VPWR VGND sg13g2_buf_8
XFILLER_97_716 VPWR VGND sg13g2_fill_1
Xfanout2620 net2625 net2620 VPWR VGND sg13g2_buf_8
XFILLER_97_749 VPWR VGND sg13g2_decap_8
Xfanout2631 net2632 net2631 VPWR VGND sg13g2_buf_8
Xfanout2642 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ net2642 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[250\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xfanout2653 net2654 net2653 VPWR VGND sg13g2_buf_8
Xfanout2697 net2698 net2697 VPWR VGND sg13g2_buf_2
XFILLER_78_952 VPWR VGND sg13g2_decap_8
Xfanout2675 net2676 net2675 VPWR VGND sg13g2_buf_8
Xfanout2664 data_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2664 VPWR
+ VGND sg13g2_buf_8
Xfanout2686 data_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2686 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] net637 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_93_944 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y
+ VPWR VGND sg13g2_nor4_1
XFILLER_65_635 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C i_snitch.pc_d\[18\]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y
+ i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C_Y VPWR
+ VGND i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B_X sg13g2_nand4_1
XFILLER_18_562 VPWR VGND sg13g2_fill_2
XFILLER_64_178 VPWR VGND sg13g2_fill_2
XFILLER_33_521 VPWR VGND sg13g2_fill_1
XFILLER_33_554 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xclkload30 clknet_leaf_44_clk clkload30/X VPWR VGND sg13g2_buf_8
Xclkload52 clknet_leaf_74_clk clkload52/X VPWR VGND sg13g2_buf_8
Xclkload41 clkload41/Y clknet_leaf_87_clk VPWR VGND sg13g2_inv_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y net2971
+ net2955 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 VPWR VGND sg13g2_nor2_2
Xclkload63 clkload63/Y clknet_leaf_82_clk VPWR VGND sg13g2_inv_2
XFILLER_88_727 VPWR VGND sg13g2_fill_2
XFILLER_96_771 VPWR VGND sg13g2_fill_1
XFILLER_84_933 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q
+ net3197 VGND VPWR net626 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_95_292 VPWR VGND sg13g2_fill_2
XFILLER_56_646 VPWR VGND sg13g2_decap_8
XFILLER_83_465 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C
+ net48 net34 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor3_2
XFILLER_70_104 VPWR VGND sg13g2_decap_4
XFILLER_55_189 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[263\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[375\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net904 net2647 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_51_340 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_fill_2
XFILLER_34_47 VPWR VGND sg13g2_decap_4
XFILLER_8_709 VPWR VGND sg13g2_fill_2
XFILLER_12_749 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ net2941 net40 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
Xclkload2 clknet_5_23__leaf_clk clkload2/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[270\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_106_843 VPWR VGND sg13g2_decap_8
XFILLER_4_948 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[376\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[376\]
+ net3137 i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
XFILLER_105_364 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y
+ net96 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
XFILLER_94_708 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C
+ net2613 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_59_99 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2
+ net2507 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_87_782 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_46_101 VPWR VGND sg13g2_fill_1
XFILLER_90_903 VPWR VGND sg13g2_decap_8
XFILLER_74_443 VPWR VGND sg13g2_fill_2
XFILLER_46_145 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[405\] clknet_leaf_114_clk sg13g2_dfrbpq_1
XFILLER_74_498 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2816 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_27_392 VPWR VGND sg13g2_fill_2
XFILLER_30_579 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR net427 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
Xhold709 i_snitch.i_snitch_regfile.mem\[128\] VPWR VGND net741 sg13g2_dlygate4sd3_1
XFILLER_10_281 VPWR VGND sg13g2_decap_4
XFILLER_7_753 VPWR VGND sg13g2_decap_8
XFILLER_7_797 VPWR VGND sg13g2_decap_8
Xfanout3140 net3140 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_buf_16
XFILLER_69_226 VPWR VGND sg13g2_fill_2
Xi_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y net1245
+ net2487 i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 VPWR VGND
+ sg13g2_nor2_1
Xfanout3162 net1404 net3162 VPWR VGND sg13g2_buf_8
Xfanout3151 i_snitch.i_snitch_lsu.metadata_q\[3\] net3151 VPWR VGND sg13g2_buf_8
Xfanout3173 i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q net3173
+ VPWR VGND sg13g2_buf_8
XFILLER_97_557 VPWR VGND sg13g2_decap_8
Xfanout3195 net3197 net3195 VPWR VGND sg13g2_buf_8
XFILLER_2_480 VPWR VGND sg13g2_fill_1
Xfanout3184 net3194 net3184 VPWR VGND sg13g2_buf_8
Xfanout2450 i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y net2450 VPWR
+ VGND sg13g2_buf_8
Xfanout2472 net2474 net2472 VPWR VGND sg13g2_buf_8
Xfanout2461 net2462 net2461 VPWR VGND sg13g2_buf_8
XFILLER_97_579 VPWR VGND sg13g2_decap_8
Xfanout2494 net2497 net2494 VPWR VGND sg13g2_buf_8
Xfanout2483 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y
+ net2483 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net883 net2680 net3041 VPWR VGND sg13g2_a22oi_1
Xrsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[111\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_81_914 VPWR VGND sg13g2_decap_8
XFILLER_66_988 VPWR VGND sg13g2_decap_4
XFILLER_66_966 VPWR VGND sg13g2_fill_2
XFILLER_80_402 VPWR VGND sg13g2_fill_2
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_19_871 VPWR VGND sg13g2_decap_4
XFILLER_19_893 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[290\] clknet_leaf_109_clk sg13g2_dfrbpq_1
XFILLER_33_373 VPWR VGND sg13g2_fill_1
XFILLER_60_170 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2548 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C
+ net2565 sg13g2_a21oi_1
XFILLER_103_802 VPWR VGND sg13g2_decap_8
XFILLER_102_301 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[425\] clknet_leaf_105_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[483\]_sg13g2_nor3_1_A net1277 net2854 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[214\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net1106 net2651 net2791 VPWR VGND sg13g2_a22oi_1
XFILLER_103_879 VPWR VGND sg13g2_decap_8
XFILLER_102_378 VPWR VGND sg13g2_decap_8
XFILLER_69_760 VPWR VGND sg13g2_fill_1
XFILLER_57_900 VPWR VGND sg13g2_fill_2
XFILLER_29_602 VPWR VGND sg13g2_fill_2
XFILLER_84_763 VPWR VGND sg13g2_fill_2
XFILLER_56_454 VPWR VGND sg13g2_decap_4
XFILLER_45_46 VPWR VGND sg13g2_fill_2
XFILLER_43_104 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\] net566 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A
+ VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND sg13g2_inv_1
XFILLER_80_980 VPWR VGND sg13g2_decap_8
XFILLER_71_479 VPWR VGND sg13g2_decap_8
XFILLER_101_63 VPWR VGND sg13g2_decap_8
XFILLER_52_682 VPWR VGND sg13g2_fill_1
XFILLER_51_170 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_12_579 VPWR VGND sg13g2_fill_1
XFILLER_40_877 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y net2846 i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1
+ net2753 net3081 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2760 net71 VPWR VGND sg13g2_nand2_1
XFILLER_106_695 VPWR VGND sg13g2_fill_2
XFILLER_106_662 VPWR VGND sg13g2_decap_8
XFILLER_105_161 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ VPWR shift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 VGND net3170 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]
+ sg13g2_o21ai_1
Xshift_reg_q\[6\]_sg13g2_nor2_1_A net506 net2731 shift_reg_q\[6\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_0_940 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[124\]
+ net2950 i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2485 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_Y net2449 net2867 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_dfrbpq_1_Q_D
+ net2912 sg13g2_a221oi_1
XFILLER_94_527 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[1\]
+ VGND i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1 net2292 sg13g2_o21ai_1
XFILLER_94_549 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B_sg13g2_nor2_1_Y
+ net2592 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2792
+ net2668 VPWR VGND sg13g2_nand2_1
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_90_799 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2490 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_37_1024 VPWR VGND sg13g2_decap_4
XFILLER_15_395 VPWR VGND sg13g2_decap_8
XFILLER_31_822 VPWR VGND sg13g2_fill_2
XFILLER_31_888 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ net2546 VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[445\] clknet_leaf_95_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[234\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net1028 net2437 net2282 VPWR VGND sg13g2_a22oi_1
Xhold517 shift_reg_q\[12\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net549 sg13g2_dlygate4sd3_1
Xshift_reg_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2728 shift_reg_q\[17\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[13\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[13\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold506 shift_reg_q\[9\] VPWR VGND net538 sg13g2_dlygate4sd3_1
Xhold528 i_snitch.sb_q\[10\] VPWR VGND net560 sg13g2_dlygate4sd3_1
Xhold539 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\] VPWR
+ VGND net571 sg13g2_dlygate4sd3_1
XFILLER_98_822 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_805 VPWR VGND sg13g2_decap_8
XFILLER_98_899 VPWR VGND sg13g2_decap_8
Xfanout2280 net2281 net2280 VPWR VGND sg13g2_buf_8
XFILLER_25_0 VPWR VGND sg13g2_decap_8
Xhold1206 i_snitch.i_snitch_regfile.mem\[194\] VPWR VGND net1238 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0 net3013 i_snitch.i_snitch_regfile.mem\[321\]
+ i_snitch.i_snitch_regfile.mem\[353\] i_snitch.i_snitch_regfile.mem\[449\] i_snitch.i_snitch_regfile.mem\[481\]
+ net2963 i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold1239 rsp_data_q\[23\] VPWR VGND net1271 sg13g2_dlygate4sd3_1
Xhold1217 i_snitch.i_snitch_regfile.mem\[485\] VPWR VGND net1249 sg13g2_dlygate4sd3_1
Xhold1228 i_snitch.i_snitch_regfile.mem\[301\] VPWR VGND net1260 sg13g2_dlygate4sd3_1
Xfanout2291 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ net2291 VPWR VGND sg13g2_buf_8
XFILLER_93_571 VPWR VGND sg13g2_fill_1
XFILLER_93_560 VPWR VGND sg13g2_decap_8
XFILLER_81_711 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR net746 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_81_755 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2886
+ net2897 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_60_clk clknet_5_31__leaf_clk clknet_leaf_60_clk VPWR VGND sg13g2_buf_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X VGND VPWR i_req_arb.gen_arbiter.req_d\[1\]
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B net1398 sg13g2_or2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 VPWR VGND i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A net763 i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B
+ i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xrsp_data_q\[26\]_sg13g2_dfrbpq_1_Q net3234 VGND VPWR rsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[26\] clknet_leaf_33_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_1 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_1_Y
+ net2983 i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_nand2b_1_A_N_Y net3009 i_snitch.i_snitch_regfile.mem\[63\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0 net3129 i_snitch.i_snitch_regfile.mem\[402\]
+ i_snitch.i_snitch_regfile.mem\[434\] i_snitch.i_snitch_regfile.mem\[466\] i_snitch.i_snitch_regfile.mem\[498\]
+ net3108 i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_103_7 VPWR VGND sg13g2_decap_8
Xoutput15 net15 uio_out[6] VPWR VGND sg13g2_buf_1
XFILLER_89_811 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y net3089
+ i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_88_343 VPWR VGND sg13g2_fill_2
XFILLER_1_748 VPWR VGND sg13g2_decap_8
XFILLER_89_888 VPWR VGND sg13g2_decap_8
XFILLER_88_354 VPWR VGND sg13g2_fill_2
XFILLER_102_175 VPWR VGND sg13g2_decap_8
XFILLER_88_387 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_and3_1_X
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A
+ i_req_arb.data_i\[39\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ net2535 VPWR VGND sg13g2_and3_1
XFILLER_29_421 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_56_251 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2442 net2771 i_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[465\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_72_788 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[254\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net921 net2437 net2244 VPWR VGND sg13g2_a22oi_1
XFILLER_32_608 VPWR VGND sg13g2_decap_4
XFILLER_72_66 VPWR VGND sg13g2_fill_1
XFILLER_13_833 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_51_clk clknet_5_26__leaf_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net1256 net2486 i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[29\]_sg13g2_nand2_1_B i_snitch.pc_d\[29\]_sg13g2_nand2_1_B_Y i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_67_1028 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1
+ VGND net2818 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_106_481 VPWR VGND sg13g2_decap_8
XFILLER_97_63 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y_sg13g2_and4_1_C
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1
+ VPWR VGND sg13g2_and4_1
XFILLER_79_332 VPWR VGND sg13g2_decap_4
XFILLER_95_814 VPWR VGND sg13g2_fill_1
XFILLER_79_365 VPWR VGND sg13g2_fill_2
XFILLER_79_354 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2444 VPWR VGND sg13g2_nand2_1
XFILLER_95_847 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A
+ VGND i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ VGND sg13g2_inv_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_or2_1_X
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D
+ net3081 net3083 sg13g2_or2_1
Xclkbuf_leaf_42_clk clknet_5_11__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1183 net2494 net1156 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0 net3122 i_snitch.i_snitch_regfile.mem\[128\]
+ i_snitch.i_snitch_regfile.mem\[160\] i_snitch.i_snitch_regfile.mem\[192\] i_snitch.i_snitch_regfile.mem\[224\]
+ net3104 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_15_181 VPWR VGND sg13g2_decap_8
XFILLER_30_140 VPWR VGND sg13g2_fill_2
XFILLER_11_1005 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ net2631 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ VPWR strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B VGND
+ net3168 net533 sg13g2_o21ai_1
XFILLER_7_94 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[99\]_sg13g2_nor3_1_A net1364 net2866 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[485\] clknet_leaf_110_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_inv_1_A_Y net3002 sg13g2_o21ai_1
XFILLER_98_685 VPWR VGND sg13g2_decap_4
Xdata_pdata\[28\]_sg13g2_nand2b_1_B data_pdata\[28\]_sg13g2_nand2b_1_B_Y data_pdata\[28\]
+ VPWR VGND net3159 sg13g2_nand2b_2
Xhold1003 data_pdata\[14\] VPWR VGND net1035 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net989 net2434 net2272 VPWR VGND sg13g2_a22oi_1
Xhold1014 i_snitch.i_snitch_regfile.mem\[45\] VPWR VGND net1046 sg13g2_dlygate4sd3_1
Xhold1058 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1090 sg13g2_dlygate4sd3_1
Xhold1036 i_snitch.i_snitch_regfile.mem\[427\] VPWR VGND net1068 sg13g2_dlygate4sd3_1
Xhold1047 i_snitch.i_snitch_regfile.mem\[43\] VPWR VGND net1079 sg13g2_dlygate4sd3_1
Xhold1025 i_snitch.i_snitch_regfile.mem\[49\] VPWR VGND net1057 sg13g2_dlygate4sd3_1
Xhold1069 i_snitch.i_snitch_regfile.mem\[422\] VPWR VGND net1101 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y net532 VPWR i_snitch.sb_d\[8\] VGND net2292 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_26_48 VPWR VGND sg13g2_fill_1
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_38_295 VPWR VGND sg13g2_fill_2
XFILLER_54_788 VPWR VGND sg13g2_fill_1
XFILLER_53_254 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_33_clk clknet_5_9__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[355\]_sg13g2_nor3_1_A net1206 net2879 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2489 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X
+ sg13g2_o21ai_1
XFILLER_22_696 VPWR VGND sg13g2_fill_1
XFILLER_42_47 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2266 net2387 net1179 VPWR VGND sg13g2_a22oi_1
XFILLER_10_847 VPWR VGND sg13g2_fill_1
XFILLER_10_858 VPWR VGND sg13g2_decap_4
Xdata_pdata\[27\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net942 data_pdata\[27\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2872
+ net2659 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q net3286 VGND VPWR i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[304\] clknet_leaf_87_clk sg13g2_dfrbpq_1
Xhold870 data_pdata\[12\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net902 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0 net3126 i_snitch.i_snitch_regfile.mem\[285\]
+ i_snitch.i_snitch_regfile.mem\[317\] i_snitch.i_snitch_regfile.mem\[349\] i_snitch.i_snitch_regfile.mem\[381\]
+ net3106 i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold881 i_snitch.i_snitch_regfile.mem\[202\] VPWR VGND net913 sg13g2_dlygate4sd3_1
XFILLER_104_963 VPWR VGND sg13g2_decap_8
Xhold892 i_snitch.i_snitch_regfile.mem\[159\] VPWR VGND net924 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B net2837
+ i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_49_505 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[67\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[67\]
+ i_snitch.i_snitch_regfile.mem\[99\] net3120 i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net505 net2324 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_92_817 VPWR VGND sg13g2_fill_2
XFILLER_92_806 VPWR VGND sg13g2_decap_8
XFILLER_76_368 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y net1174 VPWR i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A
+ VGND net2302 net2518 sg13g2_o21ai_1
XFILLER_64_508 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2380
+ sg13g2_o21ai_1
XFILLER_91_316 VPWR VGND sg13g2_decap_8
XFILLER_91_305 VPWR VGND sg13g2_fill_2
XFILLER_76_379 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_Y i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_84_390 VPWR VGND sg13g2_fill_1
XFILLER_72_541 VPWR VGND sg13g2_fill_2
XFILLER_17_435 VPWR VGND sg13g2_fill_2
XFILLER_33_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_5_3__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_12_151 VPWR VGND sg13g2_fill_1
XFILLER_40_471 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2347
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_40_493 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[294\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2899 net2779 net2317 net1209 VPWR VGND sg13g2_a22oi_1
XFILLER_4_361 VPWR VGND sg13g2_fill_2
XFILLER_4_350 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0 net3119 i_snitch.i_snitch_regfile.mem\[409\]
+ i_snitch.i_snitch_regfile.mem\[441\] i_snitch.i_snitch_regfile.mem\[473\] i_snitch.i_snitch_regfile.mem\[505\]
+ net3100 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_68_814 VPWR VGND sg13g2_fill_1
Xdata_pdata\[19\]_sg13g2_a21oi_1_A2 VGND VPWR net3158 data_pdata\[19\] data_pdata\[19\]_sg13g2_a21oi_1_A2_Y
+ net3151 sg13g2_a21oi_1
XFILLER_79_184 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y net1235 VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1 net2831
+ VPWR i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_83_828 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_B1
+ net593 net2869 VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[295\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[295\]
+ net3002 i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_a21oi_1_A1_Y net2975 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B_Y VPWR
+ VGND sg13g2_nand2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B_Y
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2662 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[429\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2381 net805 net2689 net2862 VPWR VGND sg13g2_a22oi_1
XFILLER_90_393 VPWR VGND sg13g2_fill_2
XFILLER_24_939 VPWR VGND sg13g2_fill_1
XFILLER_92_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_5_6__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_32_994 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[324\] clknet_leaf_107_clk sg13g2_dfrbpq_1
XFILLER_12_28 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[113\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2411 net922 net2664 net2870 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2610 VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1
+ VGND i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ sg13g2_o21ai_1
XFILLER_105_738 VPWR VGND sg13g2_fill_1
XFILLER_104_259 VPWR VGND sg13g2_decap_8
XFILLER_99_972 VPWR VGND sg13g2_decap_8
XFILLER_59_803 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[12\]_sg13g2_a22oi_1_A1 shift_reg_q\[12\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_mux2_1_A1_1_X
+ net3057 net3047 shift_reg_q\[12\] VPWR VGND sg13g2_a22oi_1
XFILLER_101_966 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ net2696 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_100_454 VPWR VGND sg13g2_fill_2
XFILLER_74_828 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2469
+ net2267 net2662 net2878 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VGND net2586 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_14_405 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]
+ net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2465
+ net2274 net2687 net2862 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1
+ net1396 VGND sg13g2_inv_1
XFILLER_41_279 VPWR VGND sg13g2_fill_2
XFILLER_22_493 VPWR VGND sg13g2_fill_2
XFILLER_6_615 VPWR VGND sg13g2_fill_1
XFILLER_6_604 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_B
+ net98 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y
+ sg13g2_nand4_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.inst_addr_o\[31\] net2524 VPWR VGND sg13g2_xnor2_1
XFILLER_5_158 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2543 VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_2_810 VPWR VGND sg13g2_decap_8
Xfanout2802 net2809 net2802 VPWR VGND sg13g2_buf_8
Xfanout2835 i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1_B1 net2835 VPWR
+ VGND sg13g2_buf_8
Xfanout2824 net2825 net2824 VPWR VGND sg13g2_buf_8
Xfanout2813 i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1_A2 net2813 VPWR
+ VGND sg13g2_buf_8
Xfanout2846 net2847 net2846 VPWR VGND sg13g2_buf_8
XFILLER_89_482 VPWR VGND sg13g2_fill_1
Xfanout2857 net2859 net2857 VPWR VGND sg13g2_buf_8
XFILLER_49_324 VPWR VGND sg13g2_fill_1
XFILLER_2_887 VPWR VGND sg13g2_decap_8
Xfanout2868 net2869 net2868 VPWR VGND sg13g2_buf_8
Xfanout2879 net2880 net2879 VPWR VGND sg13g2_buf_8
XFILLER_94_42 VPWR VGND sg13g2_decap_8
XFILLER_76_154 VPWR VGND sg13g2_decap_8
XFILLER_64_349 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_dfrbpq_1_Q net3315 VGND VPWR i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[344\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_A1
+ net2309 i_snitch.pc_d\[14\] i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
XFILLER_72_360 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_21_909 VPWR VGND sg13g2_fill_1
XFILLER_14_983 VPWR VGND sg13g2_fill_1
Xi_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q net3251 VGND VPWR i_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.gpr_waddr\[6\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_43_90 VPWR VGND sg13g2_fill_2
XFILLER_9_453 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3091 i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
Xuio_out_sg13g2_inv_1_Y VPWR net12 uio_out_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_4_84 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_4_clk clknet_5_4__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
XFILLER_96_964 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ net2716 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_83_636 VPWR VGND sg13g2_decap_8
XFILLER_55_338 VPWR VGND sg13g2_decap_4
XFILLER_71_809 VPWR VGND sg13g2_fill_1
XFILLER_64_883 VPWR VGND sg13g2_decap_8
XFILLER_17_1000 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2347
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] VGND sg13g2_inv_1
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_32_791 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VGND sg13g2_inv_1
XFILLER_20_975 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[469\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net943 net2460 net2268 VPWR VGND sg13g2_a22oi_1
Xshift_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2730 shift_reg_q\[5\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[1\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y net3001 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2364
+ sg13g2_o21ai_1
Xuo_out_sg13g2_buf_1_X_5 i_req_register.data_o\[39\] net22 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y
+ net3175 net1319 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[364\] clknet_leaf_70_clk sg13g2_dfrbpq_1
XFILLER_63_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net1151 net2445 net2266 VPWR VGND sg13g2_a22oi_1
XFILLER_48_35 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[227\]_sg13g2_nor3_1_A net1327 net2873 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_100_240 VPWR VGND sg13g2_decap_8
XFILLER_87_986 VPWR VGND sg13g2_decap_8
XFILLER_104_63 VPWR VGND sg13g2_decap_8
XFILLER_73_102 VPWR VGND sg13g2_fill_2
XFILLER_46_338 VPWR VGND sg13g2_fill_1
XFILLER_73_157 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[384\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand4_1_Y
+ net2925 net2922 net3033 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.inst_addr_o\[23\] net2526 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ net3007 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_nor3_1
XFILLER_55_883 VPWR VGND sg13g2_fill_1
XFILLER_42_522 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[490\]
+ net2801 i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xdata_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A
+ data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ VGND sg13g2_inv_2
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1_sg13g2_and2_1_X i_snitch.inst_addr_o\[17\]
+ net2528 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1 VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]
+ net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_6_412 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[24\]_sg13g2_dfrbpq_1_Q net3313 VGND VPWR i_snitch.pc_d\[24\]
+ i_snitch.inst_addr_o\[24\] clknet_leaf_54_clk sg13g2_dfrbpq_2
Xfanout3322 net3324 net3322 VPWR VGND sg13g2_buf_8
Xfanout3311 net3313 net3311 VPWR VGND sg13g2_buf_8
Xfanout3300 net3301 net3300 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2574 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xfanout2610 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X
+ net2610 VPWR VGND sg13g2_buf_8
Xfanout2621 net2625 net2621 VPWR VGND sg13g2_buf_8
Xfanout2632 net2633 net2632 VPWR VGND sg13g2_buf_8
Xfanout2643 data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ net2643 VPWR VGND sg13g2_buf_8
XFILLER_2_684 VPWR VGND sg13g2_decap_8
Xfanout2654 data_pdata\[29\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2654 VPWR
+ VGND sg13g2_buf_8
Xrsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_77_441 VPWR VGND sg13g2_fill_1
Xfanout2665 net2666 net2665 VPWR VGND sg13g2_buf_8
Xfanout2676 data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2676 VPWR VGND sg13g2_buf_8
Xfanout2687 data_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2687 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2594 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_nand2_1
Xfanout2698 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ net2698 VPWR VGND sg13g2_buf_8
XFILLER_93_923 VPWR VGND sg13g2_decap_8
XFILLER_92_400 VPWR VGND sg13g2_decap_8
XFILLER_65_603 VPWR VGND sg13g2_fill_1
XFILLER_64_168 VPWR VGND sg13g2_fill_1
XFILLER_18_596 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[489\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2367 net875 net2685 net2855 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net123 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
XFILLER_14_791 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[384\] clknet_leaf_18_clk sg13g2_dfrbpq_1
Xclkload20 clknet_leaf_38_clk clkload20/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[173\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2344 net1002 net2690 net2774 VPWR VGND sg13g2_a22oi_1
Xclkload31 clknet_leaf_45_clk clkload31/Y VPWR VGND sg13g2_inv_4
Xclkload53 clknet_leaf_52_clk clkload53/X VPWR VGND sg13g2_buf_8
Xclkload42 clkload42/Y clknet_leaf_89_clk VPWR VGND sg13g2_inv_2
Xclkload64 clkload64/Y clknet_leaf_55_clk VPWR VGND sg13g2_inv_8
XFILLER_88_706 VPWR VGND sg13g2_decap_8
XFILLER_69_920 VPWR VGND sg13g2_fill_2
XFILLER_96_750 VPWR VGND sg13g2_decap_8
XFILLER_68_430 VPWR VGND sg13g2_fill_1
XFILLER_84_912 VPWR VGND sg13g2_decap_8
XFILLER_68_452 VPWR VGND sg13g2_decap_4
XFILLER_83_433 VPWR VGND sg13g2_decap_4
XFILLER_68_496 VPWR VGND sg13g2_fill_2
XFILLER_18_27 VPWR VGND sg13g2_fill_1
XFILLER_84_989 VPWR VGND sg13g2_decap_8
XFILLER_83_455 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2629 net2851 net74
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2672 net2780 net2318 net1195 VPWR VGND sg13g2_a22oi_1
XFILLER_43_319 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_24_555 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B_sg13g2_or4_1_X
+ net3146 net109 net3085 net3087 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_or4_1
XFILLER_52_897 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[203\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xclkload3 clknet_5_27__leaf_clk clkload3/X VPWR VGND sg13g2_buf_8
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\] net2622 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_106_822 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[309\]
+ net3005 i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_a21oi_1_A1_Y net2978 sg13g2_a21oi_1
XFILLER_4_927 VPWR VGND sg13g2_decap_8
XFILLER_105_343 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y net2933 sg13g2_a21oi_2
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y net491 VPWR i_snitch.sb_d\[15\] VGND net2292
+ i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_3_437 VPWR VGND sg13g2_fill_2
XFILLER_106_899 VPWR VGND sg13g2_decap_8
XFILLER_79_728 VPWR VGND sg13g2_fill_1
XFILLER_59_56 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ VPWR VGND sg13g2_nand2_2
Xcnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net543 cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 VPWR VGND sg13g2_nand2_1
XFILLER_75_901 VPWR VGND sg13g2_fill_1
XFILLER_74_422 VPWR VGND sg13g2_decap_4
XFILLER_74_411 VPWR VGND sg13g2_fill_2
XFILLER_90_959 VPWR VGND sg13g2_decap_8
XFILLER_15_500 VPWR VGND sg13g2_decap_4
XFILLER_91_32 VPWR VGND sg13g2_fill_1
XFILLER_91_21 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ net3087 net122 VPWR VGND sg13g2_nand2_2
XFILLER_61_138 VPWR VGND sg13g2_decap_8
XFILLER_43_853 VPWR VGND sg13g2_fill_1
XFILLER_43_842 VPWR VGND sg13g2_fill_2
XFILLER_43_831 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1
+ VGND net2610 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A
+ sg13g2_o21ai_1
XFILLER_11_772 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2360 net841 net2685 net2767 VPWR VGND sg13g2_a22oi_1
XFILLER_7_776 VPWR VGND sg13g2_fill_1
Xfanout3130 net3131 net3130 VPWR VGND sg13g2_buf_8
Xfanout3141 net109 net3141 VPWR VGND sg13g2_buf_8
Xfanout3174 net3176 net3174 VPWR VGND sg13g2_buf_8
Xfanout3152 net3153 net3152 VPWR VGND sg13g2_buf_8
Xfanout3163 net1402 net3163 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_a22oi_1_B2_Y
+ net2403 net664 net2644 net2796 VPWR VGND sg13g2_a22oi_1
Xfanout3196 net3197 net3196 VPWR VGND sg13g2_buf_8
Xfanout2451 net2452 net2451 VPWR VGND sg13g2_buf_8
Xfanout3185 net3194 net3185 VPWR VGND sg13g2_buf_8
Xfanout2440 net2441 net2440 VPWR VGND sg13g2_buf_8
Xfanout2462 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2462 VPWR
+ VGND sg13g2_buf_8
Xfanout2495 net2497 net2495 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]
+ net3170 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_27_4 VPWR VGND sg13g2_decap_8
Xfanout2484 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2484 VPWR VGND sg13g2_buf_8
Xfanout2473 net2474 net2473 VPWR VGND sg13g2_buf_8
XFILLER_93_742 VPWR VGND sg13g2_decap_4
XFILLER_78_783 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[42\]
+ net2827 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_a21oi_1_A1_Y net2822 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_nor3_1_A net1286 net2885 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q net3305 VGND VPWR i_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[223\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2959
+ i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2965
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_77_1019 VPWR VGND sg13g2_decap_8
XFILLER_65_499 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[4\]_sg13g2_nor2_1_A net472 net2727 strb_reg_q\[4\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A
+ VGND net2540 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.gpr_waddr\[7\]_sg13g2_nand2_1_A data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D
+ i_snitch.gpr_waddr\[7\] i_snitch.gpr_waddr\[6\] VPWR VGND sg13g2_nand2_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1
+ net712 net622 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_A_N i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_B1
+ i_snitch.inst_addr_o\[14\] i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1 VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ net2684 net2745 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_88_503 VPWR VGND sg13g2_fill_1
XFILLER_0_407 VPWR VGND sg13g2_decap_8
XFILLER_103_858 VPWR VGND sg13g2_decap_8
XFILLER_102_357 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1
+ sg13g2_a21oi_1
XFILLER_96_580 VPWR VGND sg13g2_fill_2
XFILLER_56_422 VPWR VGND sg13g2_fill_2
Xdata_pdata\[11\]_sg13g2_nor2b_1_A data_pdata\[11\] net3158 data_pdata\[11\]_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_84_753 VPWR VGND sg13g2_fill_1
XFILLER_84_742 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_83_296 VPWR VGND sg13g2_fill_2
XFILLER_101_42 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2360 net923 net2456 net2251 VPWR VGND sg13g2_a22oi_1
XFILLER_24_396 VPWR VGND sg13g2_fill_1
XFILLER_25_897 VPWR VGND sg13g2_fill_1
XFILLER_61_46 VPWR VGND sg13g2_decap_4
XFILLER_8_507 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ net2589 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_61_79 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[348\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net909 net2473 net2246 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[243\] clknet_leaf_121_clk sg13g2_dfrbpq_1
XFILLER_3_212 VPWR VGND sg13g2_decap_8
XFILLER_105_140 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_fill_1
XFILLER_86_54 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y
+ net2642 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A
+ VPWR VGND sg13g2_nor3_1
XFILLER_102_891 VPWR VGND sg13g2_decap_8
XFILLER_75_720 VPWR VGND sg13g2_decap_4
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B_sg13g2_and2_1_X
+ i_snitch.inst_addr_o\[19\] net2525 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_and2_1
XFILLER_0_996 VPWR VGND sg13g2_decap_8
XFILLER_74_230 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[7\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR rsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[7\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_16_853 VPWR VGND sg13g2_fill_1
XFILLER_15_352 VPWR VGND sg13g2_fill_1
XFILLER_96_7 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[9\] net991 net2914 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_30_366 VPWR VGND sg13g2_decap_4
Xhold518 shift_reg_q\[26\] VPWR VGND net550 sg13g2_dlygate4sd3_1
Xhold507 shift_reg_q\[9\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net539 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\] net660 net2620
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xhold529 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\] VPWR
+ VGND net561 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B
+ net2959 i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_98_801 VPWR VGND sg13g2_decap_8
XFILLER_83_1012 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_97_344 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2428 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_98_878 VPWR VGND sg13g2_decap_8
XFILLER_97_377 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q
+ net3230 VGND VPWR net595 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_1
Xfanout2270 net2271 net2270 VPWR VGND sg13g2_buf_8
Xhold1207 i_snitch.i_snitch_regfile.mem\[165\] VPWR VGND net1239 sg13g2_dlygate4sd3_1
XFILLER_97_388 VPWR VGND sg13g2_decap_8
Xfanout2281 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B_X
+ net2281 VPWR VGND sg13g2_buf_8
Xfanout2292 net2293 net2292 VPWR VGND sg13g2_buf_8
Xhold1229 i_snitch.i_snitch_regfile.mem\[498\] VPWR VGND net1261 sg13g2_dlygate4sd3_1
Xhold1218 i_snitch.i_snitch_regfile.mem\[122\] VPWR VGND net1250 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[81\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2355 net1203 net2664 net2786 VPWR VGND sg13g2_a22oi_1
XFILLER_39_934 VPWR VGND sg13g2_fill_1
XFILLER_39_967 VPWR VGND sg13g2_decap_4
XFILLER_66_775 VPWR VGND sg13g2_fill_1
XFILLER_38_466 VPWR VGND sg13g2_fill_2
XFILLER_53_436 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net1094 net2470 net2263 VPWR VGND sg13g2_a22oi_1
XFILLER_53_469 VPWR VGND sg13g2_decap_4
XFILLER_22_812 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1
+ VPWR VGND net3142 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[263\] clknet_leaf_118_clk sg13g2_dfrbpq_1
XFILLER_21_355 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q
+ net3245 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[407\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[369\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[369\]
+ net3135 i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
XFILLER_1_727 VPWR VGND sg13g2_decap_8
Xoutput16 net16 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_103_644 VPWR VGND sg13g2_decap_8
XFILLER_103_622 VPWR VGND sg13g2_fill_1
XFILLER_89_867 VPWR VGND sg13g2_decap_8
XFILLER_0_237 VPWR VGND sg13g2_fill_1
XFILLER_103_655 VPWR VGND sg13g2_fill_1
XFILLER_102_154 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[389\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_57_731 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2417 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_5_1012 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[259\] net2814 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ net2631 VPWR i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
XFILLER_56_230 VPWR VGND sg13g2_fill_2
XFILLER_45_904 VPWR VGND sg13g2_fill_1
XFILLER_84_550 VPWR VGND sg13g2_fill_2
XFILLER_71_200 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3172 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ state sg13g2_a21oi_1
XFILLER_56_263 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2701 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_17_639 VPWR VGND sg13g2_fill_2
XFILLER_72_778 VPWR VGND sg13g2_decap_8
XFILLER_71_255 VPWR VGND sg13g2_fill_1
XFILLER_71_244 VPWR VGND sg13g2_decap_4
XFILLER_60_929 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2_sg13g2_and3_1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_and3_1
XFILLER_25_683 VPWR VGND sg13g2_fill_1
XFILLER_40_642 VPWR VGND sg13g2_fill_1
XFILLER_8_315 VPWR VGND sg13g2_fill_1
XFILLER_12_377 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2442 net2771 i_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR net567 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ net2607 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B net2867 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_2
XFILLER_97_42 VPWR VGND sg13g2_decap_8
XFILLER_67_506 VPWR VGND sg13g2_fill_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B_sg13g2_o21ai_1_Y
+ net2525 VPWR i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B
+ VGND i_snitch.inst_addr_o\[19\] i_snitch.inst_addr_o\[20\] sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C
+ net3034 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A
+ net2922 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B
+ VPWR VGND sg13g2_and4_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_0_793 VPWR VGND sg13g2_decap_8
XFILLER_11_7 VPWR VGND sg13g2_decap_8
XFILLER_75_572 VPWR VGND sg13g2_decap_8
XFILLER_75_561 VPWR VGND sg13g2_fill_1
XFILLER_75_550 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_47_263 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[283\] clknet_leaf_119_clk sg13g2_dfrbpq_1
XFILLER_75_594 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2707 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_50_439 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VGND net2702 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2641 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[418\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[418\] clknet_leaf_13_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[207\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2339 net1080 net2678 net2793 VPWR VGND sg13g2_a22oi_1
XFILLER_98_653 VPWR VGND sg13g2_decap_4
XFILLER_86_804 VPWR VGND sg13g2_fill_1
XFILLER_58_506 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y net3089
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y sg13g2_o21ai_1
Xhold1004 data_pdata\[14\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net1036 sg13g2_dlygate4sd3_1
Xhold1015 i_snitch.i_snitch_regfile.mem\[144\] VPWR VGND net1047 sg13g2_dlygate4sd3_1
XFILLER_100_658 VPWR VGND sg13g2_fill_2
XFILLER_100_647 VPWR VGND sg13g2_fill_1
Xhold1037 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]
+ VPWR VGND net1069 sg13g2_dlygate4sd3_1
Xhold1048 i_snitch.i_snitch_regfile.mem\[207\] VPWR VGND net1080 sg13g2_dlygate4sd3_1
Xhold1026 i_snitch.i_snitch_regfile.mem\[240\] VPWR VGND net1058 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q net3280 VGND VPWR i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[102\] clknet_leaf_76_clk sg13g2_dfrbpq_1
XFILLER_66_572 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2450 VPWR VGND sg13g2_nand2_1
Xhold1059 i_snitch.i_snitch_regfile.mem\[78\] VPWR VGND net1091 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_929 VPWR VGND sg13g2_fill_1
XFILLER_10_804 VPWR VGND sg13g2_decap_4
XFILLER_22_686 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2440 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A VPWR
+ VGND sg13g2_and2_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2 VPWR
+ VGND net2759 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_C1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2851 sg13g2_a221oi_1
XFILLER_104_942 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A
+ net3086 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xhold882 rsp_state_q VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold871 i_snitch.i_snitch_regfile.mem\[246\] VPWR VGND net903 sg13g2_dlygate4sd3_1
Xhold860 i_snitch.i_snitch_regfile.mem\[459\] VPWR VGND net892 sg13g2_dlygate4sd3_1
Xstrb_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2727 strb_reg_q\[3\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D strb_reg_q\[2\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2695 net2556 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_89_664 VPWR VGND sg13g2_decap_8
Xhold893 data_pdata\[20\] VPWR VGND net925 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0 net3007 i_snitch.i_snitch_regfile.mem\[132\]
+ i_snitch.i_snitch_regfile.mem\[164\] i_snitch.i_snitch_regfile.mem\[196\] i_snitch.i_snitch_regfile.mem\[228\]
+ net2980 i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2578 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_76_314 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y
+ net44 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2380
+ sg13g2_o21ai_1
Xshift_reg_q\[9\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net539 shift_reg_q\[9\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
XFILLER_103_496 VPWR VGND sg13g2_fill_2
XFILLER_18_904 VPWR VGND sg13g2_fill_1
XFILLER_85_892 VPWR VGND sg13g2_decap_8
XFILLER_72_520 VPWR VGND sg13g2_decap_4
XFILLER_44_255 VPWR VGND sg13g2_fill_1
XFILLER_17_447 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_Y
+ VPWR VGND i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ sg13g2_nand2b_2
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1
+ net2724 net3022 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_73_1022 VPWR VGND sg13g2_decap_8
XFILLER_72_597 VPWR VGND sg13g2_decap_4
XFILLER_26_970 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_93 VPWR VGND sg13g2_fill_1
XFILLER_41_962 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[438\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_9_635 VPWR VGND sg13g2_decap_4
XFILLER_9_624 VPWR VGND sg13g2_fill_2
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_156 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_B1
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ net2699 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C
+ net2612 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D_sg13g2_and2_1_X
+ net2569 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1 net3019 i_snitch.i_snitch_regfile.mem\[140\]
+ i_snitch.i_snitch_regfile.mem\[172\] i_snitch.i_snitch_regfile.mem\[204\] i_snitch.i_snitch_regfile.mem\[236\]
+ net2990 i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_99_417 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[122\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_a221oi_1_A1 VPWR VGND i_snitch.i_snitch_regfile.mem\[161\]
+ net3027 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[33\]
+ i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_a221oi_1_A1_Y net2831 sg13g2_a221oi_1
XFILLER_80_1015 VPWR VGND sg13g2_decap_8
XFILLER_79_130 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2422 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_83_807 VPWR VGND sg13g2_fill_1
Xi_req_arb.data_i\[41\]_sg13g2_dfrbpq_1_Q net3257 VGND VPWR i_snitch.pc_d\[6\] i_req_arb.data_i\[41\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_2
XFILLER_0_590 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2530 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2479 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[15\]_sg13g2_a21o_1_A2 i_snitch.pc_d\[15\] i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1
+ i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_B1 i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_X VPWR
+ VGND sg13g2_a21o_1
XFILLER_48_572 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2437 VPWR VGND sg13g2_nand2_1
XFILLER_36_701 VPWR VGND sg13g2_decap_4
XFILLER_48_583 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[21\]_sg13g2_dfrbpq_1_Q net3187 VGND VPWR net484 shift_reg_q\[21\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
XFILLER_90_350 VPWR VGND sg13g2_decap_8
XFILLER_91_884 VPWR VGND sg13g2_decap_8
XFILLER_51_737 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_fill_2
XFILLER_50_247 VPWR VGND sg13g2_decap_8
XFILLER_85_0 VPWR VGND sg13g2_decap_4
XFILLER_31_483 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[19\]_sg13g2_dfrbpq_1_Q net3232 VGND VPWR rsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[19\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_104_238 VPWR VGND sg13g2_decap_8
XFILLER_99_951 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net833 net702 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2638 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_85_100 VPWR VGND sg13g2_fill_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1_X
+ VPWR VGND sg13g2_and2_1
XFILLER_101_945 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1382 net2491 net1210 VPWR VGND sg13g2_a22oi_1
XFILLER_100_477 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q net3274 VGND VPWR i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[458\] clknet_leaf_103_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y
+ net109 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2761 net2308
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2519 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_54_520 VPWR VGND sg13g2_decap_4
XFILLER_26_211 VPWR VGND sg13g2_fill_1
XFILLER_27_723 VPWR VGND sg13g2_decap_4
XFILLER_39_594 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[247\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net1005 net2648 net2875 VPWR VGND sg13g2_a22oi_1
XFILLER_66_391 VPWR VGND sg13g2_fill_2
XFILLER_57_1017 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_82_895 VPWR VGND sg13g2_decap_8
XFILLER_81_372 VPWR VGND sg13g2_fill_1
XFILLER_57_1028 VPWR VGND sg13g2_fill_1
XFILLER_23_940 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1 net3018 i_snitch.i_snitch_regfile.mem\[142\]
+ i_snitch.i_snitch_regfile.mem\[174\] i_snitch.i_snitch_regfile.mem\[206\] i_snitch.i_snitch_regfile.mem\[238\]
+ net2989 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_26_299 VPWR VGND sg13g2_decap_8
XFILLER_42_748 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q net3289 VGND VPWR i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[142\] clknet_leaf_88_clk sg13g2_dfrbpq_1
XFILLER_23_984 VPWR VGND sg13g2_fill_1
XFILLER_10_623 VPWR VGND sg13g2_fill_2
Xdata_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A
+ data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ VGND sg13g2_inv_2
XFILLER_5_137 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2459 net2854 i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
Xdata_pdata\[3\]_sg13g2_nor2_1_B net3157 data_pdata\[3\] data_pdata\[3\]_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xfanout2803 net2809 net2803 VPWR VGND sg13g2_buf_2
Xhold690 data_pdata\[23\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net722 sg13g2_dlygate4sd3_1
Xfanout2814 i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2 net2814 VPWR
+ VGND sg13g2_buf_8
XFILLER_2_866 VPWR VGND sg13g2_decap_8
Xfanout2836 net2837 net2836 VPWR VGND sg13g2_buf_8
Xfanout2825 net2826 net2825 VPWR VGND sg13g2_buf_8
XFILLER_49_314 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2322
+ sg13g2_o21ai_1
Xfanout2847 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y
+ net2847 VPWR VGND sg13g2_buf_8
Xfanout2858 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y
+ net2858 VPWR VGND sg13g2_buf_8
Xfanout2869 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X net2869
+ VPWR VGND sg13g2_buf_8
XFILLER_76_122 VPWR VGND sg13g2_fill_2
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_94_21 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ net1272 VGND sg13g2_inv_1
XFILLER_64_306 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y net3088
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_92_648 VPWR VGND sg13g2_decap_8
XFILLER_76_199 VPWR VGND sg13g2_decap_4
XFILLER_64_339 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[452\]_sg13g2_nor3_1_A net1281 net2739 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_73_895 VPWR VGND sg13g2_fill_1
XFILLER_18_789 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2334
+ sg13g2_o21ai_1
XFILLER_17_299 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2603 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2365
+ sg13g2_o21ai_1
XFILLER_9_443 VPWR VGND sg13g2_decap_4
XFILLER_9_432 VPWR VGND sg13g2_fill_2
XFILLER_9_476 VPWR VGND sg13g2_decap_8
XFILLER_9_487 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2464
+ net2513 net2901 net2862 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[478\] clknet_leaf_93_clk sg13g2_dfrbpq_1
XFILLER_5_693 VPWR VGND sg13g2_fill_1
XFILLER_102_709 VPWR VGND sg13g2_decap_8
XFILLER_99_269 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2612 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2325 net787 net2680 net2893 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2379
+ sg13g2_o21ai_1
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_96_943 VPWR VGND sg13g2_decap_8
XFILLER_83_615 VPWR VGND sg13g2_decap_8
XFILLER_67_166 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0 net3136 i_snitch.i_snitch_regfile.mem\[139\]
+ i_snitch.i_snitch_regfile.mem\[171\] i_snitch.i_snitch_regfile.mem\[203\] i_snitch.i_snitch_regfile.mem\[235\]
+ net3112 i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1 net3016 i_snitch.i_snitch_regfile.mem\[144\]
+ i_snitch.i_snitch_regfile.mem\[176\] i_snitch.i_snitch_regfile.mem\[208\] i_snitch.i_snitch_regfile.mem\[240\]
+ net2987 i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2476 net2433 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2417 sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[162\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_82_158 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C_sg13g2_nand3_1_Y
+ net3077 net2927 net3083 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C
+ VPWR VGND sg13g2_nand3_1
XFILLER_51_501 VPWR VGND sg13g2_decap_4
XFILLER_90_180 VPWR VGND sg13g2_decap_4
XFILLER_63_394 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[268\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[268\]
+ net3029 i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_a21oi_1_A1_Y net2991 sg13g2_a21oi_1
XFILLER_51_567 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1 net3019 i_snitch.i_snitch_regfile.mem\[392\]
+ i_snitch.i_snitch_regfile.mem\[424\] i_snitch.i_snitch_regfile.mem\[456\] i_snitch.i_snitch_regfile.mem\[488\]
+ net2990 i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_104_1026 VPWR VGND sg13g2_fill_2
Xuo_out_sg13g2_buf_1_X_6 i_req_register.data_o\[40\] net23 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B
+ net2959 i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2413
+ sg13g2_o21ai_1
XFILLER_48_25 VPWR VGND sg13g2_fill_1
XFILLER_98_280 VPWR VGND sg13g2_fill_2
XFILLER_87_965 VPWR VGND sg13g2_decap_8
XFILLER_59_645 VPWR VGND sg13g2_fill_2
XFILLER_101_753 VPWR VGND sg13g2_decap_4
XFILLER_74_615 VPWR VGND sg13g2_decap_4
XFILLER_59_689 VPWR VGND sg13g2_decap_8
XFILLER_58_166 VPWR VGND sg13g2_decap_8
XFILLER_104_42 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2 VGND
+ VPWR net2964 i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_100_296 VPWR VGND sg13g2_decap_8
XFILLER_15_759 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2399
+ sg13g2_o21ai_1
XFILLER_70_1025 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[498\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_23_792 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[78\]
+ i_snitch.i_snitch_regfile.mem\[110\] net3130 i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_453 VPWR VGND sg13g2_fill_2
XFILLER_10_442 VPWR VGND sg13g2_fill_1
XFILLER_11_954 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2326 net917 net2645 net2894 VPWR VGND sg13g2_a22oi_1
XFILLER_10_464 VPWR VGND sg13g2_decap_4
Xfanout3312 net3313 net3312 VPWR VGND sg13g2_buf_8
Xfanout3323 net3324 net3323 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[182\] clknet_leaf_61_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1 net3016 i_snitch.i_snitch_regfile.mem\[146\]
+ i_snitch.i_snitch_regfile.mem\[178\] i_snitch.i_snitch_regfile.mem\[210\] i_snitch.i_snitch_regfile.mem\[242\]
+ net2987 i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xfanout3301 net3329 net3301 VPWR VGND sg13g2_buf_8
Xfanout2600 net2602 net2600 VPWR VGND sg13g2_buf_8
Xfanout2611 net2612 net2611 VPWR VGND sg13g2_buf_8
Xfanout2633 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y
+ net2633 VPWR VGND sg13g2_buf_8
Xfanout2644 data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ net2644 VPWR VGND sg13g2_buf_8
Xfanout2622 net2625 net2622 VPWR VGND sg13g2_buf_8
XFILLER_1_151 VPWR VGND sg13g2_fill_2
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_2_663 VPWR VGND sg13g2_decap_8
Xfanout2666 data_pdata\[24\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2666 VPWR
+ VGND sg13g2_buf_8
Xfanout2677 data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ net2677 VPWR VGND sg13g2_buf_8
Xfanout2655 net2656 net2655 VPWR VGND sg13g2_buf_8
XFILLER_29_8 VPWR VGND sg13g2_fill_1
Xfanout2688 data_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2688 VPWR VGND sg13g2_buf_8
Xfanout2699 net2703 net2699 VPWR VGND sg13g2_buf_8
XFILLER_93_902 VPWR VGND sg13g2_decap_8
XFILLER_78_987 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[106\]
+ net2953 i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_37_328 VPWR VGND sg13g2_fill_2
XFILLER_93_979 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_73_670 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y net2512
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_60_320 VPWR VGND sg13g2_fill_2
XFILLER_33_545 VPWR VGND sg13g2_decap_8
XFILLER_61_898 VPWR VGND sg13g2_fill_2
XFILLER_61_887 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[317\] clknet_leaf_95_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2854
+ net2897 VPWR VGND sg13g2_nand2_1
XFILLER_60_375 VPWR VGND sg13g2_fill_2
XFILLER_14_781 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y net2282 net2411 net1302
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1 i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A
+ i_req_arb.data_i\[39\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C net2642
+ i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y
+ VPWR VGND sg13g2_nor4_1
XFILLER_13_291 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y VPWR VGND sg13g2_and3_1
Xi_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xstrb_reg_q\[0\]_sg13g2_dfrbpq_1_Q net3184 VGND VPWR net502 strb_reg_q\[0\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
Xclkload10 clknet_leaf_4_clk clkload10/X VPWR VGND sg13g2_buf_8
Xclkload21 clknet_leaf_34_clk clkload21/X VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xclkload32 clknet_leaf_98_clk clkload32/X VPWR VGND sg13g2_buf_8
Xclkload43 clkload43/Y clknet_leaf_90_clk VPWR VGND sg13g2_inv_2
XFILLER_86_1021 VPWR VGND sg13g2_decap_8
Xclkload54 clkload54/Y clknet_leaf_53_clk VPWR VGND sg13g2_inv_2
Xclkload65 clkload65/Y clknet_leaf_67_clk VPWR VGND sg13g2_inv_2
XFILLER_6_991 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_fill_2
XFILLER_102_528 VPWR VGND sg13g2_fill_2
XFILLER_88_729 VPWR VGND sg13g2_fill_1
XFILLER_102_539 VPWR VGND sg13g2_decap_8
XFILLER_68_464 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0_X
+ net2937 net2931 i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_96_795 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2783
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_95_294 VPWR VGND sg13g2_fill_1
XFILLER_84_968 VPWR VGND sg13g2_decap_8
XFILLER_71_607 VPWR VGND sg13g2_fill_1
XFILLER_37_851 VPWR VGND sg13g2_fill_2
XFILLER_93_1014 VPWR VGND sg13g2_decap_8
XFILLER_92_990 VPWR VGND sg13g2_decap_8
XFILLER_63_180 VPWR VGND sg13g2_decap_4
XFILLER_52_854 VPWR VGND sg13g2_fill_2
XFILLER_24_534 VPWR VGND sg13g2_fill_2
XFILLER_36_394 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1 net3022 i_snitch.i_snitch_regfile.mem\[148\]
+ i_snitch.i_snitch_regfile.mem\[180\] i_snitch.i_snitch_regfile.mem\[212\] i_snitch.i_snitch_regfile.mem\[244\]
+ net2993 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y
+ i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_Y i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C_Y VPWR VGND i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_Y
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_nand2_1_A_1 i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_nand2_1_A_1_Y
+ i_snitch.i_snitch_regfile.mem\[33\] net2825 VPWR VGND sg13g2_nand2_1
Xclkload4 clknet_5_31__leaf_clk clkload4/X VPWR VGND sg13g2_buf_8
XFILLER_20_784 VPWR VGND sg13g2_fill_1
XFILLER_106_801 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2501 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ net2483 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1 net3024 i_snitch.i_snitch_regfile.mem\[396\]
+ i_snitch.i_snitch_regfile.mem\[428\] i_snitch.i_snitch_regfile.mem\[460\] i_snitch.i_snitch_regfile.mem\[492\]
+ net2991 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[29\]_sg13g2_nand2b_1_B_Y net3150 data_pdata\[21\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[13\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
XFILLER_105_322 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q net3286 VGND VPWR i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[50\] clknet_leaf_87_clk sg13g2_dfrbpq_1
XFILLER_106_878 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VGND net2599 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ sg13g2_o21ai_1
XFILLER_105_399 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[119\]
+ net2806 i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_93_209 VPWR VGND sg13g2_decap_4
XFILLER_87_762 VPWR VGND sg13g2_fill_2
XFILLER_87_795 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[504\]_sg13g2_o21ai_1_A1 net2966 VPWR i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[504\] net2806 sg13g2_o21ai_1
XFILLER_47_648 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[337\] clknet_leaf_80_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_47_659 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2450 net2245 net2411 net1216 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nor3_1_A net1237 net2784 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
XFILLER_90_938 VPWR VGND sg13g2_decap_8
XFILLER_74_478 VPWR VGND sg13g2_fill_2
XFILLER_34_309 VPWR VGND sg13g2_decap_4
XFILLER_70_640 VPWR VGND sg13g2_fill_1
XFILLER_55_692 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ net2554 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_578 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_o21ai_1_A1 net3017 VPWR i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[46\] net2988 sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B
+ VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A
+ sg13g2_or2_1
XFILLER_10_250 VPWR VGND sg13g2_fill_2
XFILLER_7_711 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[25\]_sg13g2_a22oi_1_A1 shift_reg_q\[25\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_1_X
+ net3053 net3044 shift_reg_q\[25\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y net2918 i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_6_243 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
Xfanout3120 net3121 net3120 VPWR VGND sg13g2_buf_8
Xfanout3131 net3132 net3131 VPWR VGND sg13g2_buf_8
Xfanout3142 net3143 net3142 VPWR VGND sg13g2_buf_8
Xfanout3153 net3154 net3153 VPWR VGND sg13g2_buf_8
XFILLER_3_983 VPWR VGND sg13g2_decap_8
Xfanout3164 net3165 net3164 VPWR VGND sg13g2_buf_8
Xfanout3175 net3176 net3175 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_A1
+ net2305 i_snitch.pc_d\[25\] i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xfanout3197 net3205 net3197 VPWR VGND sg13g2_buf_8
XFILLER_2_460 VPWR VGND sg13g2_decap_4
Xfanout3186 net3188 net3186 VPWR VGND sg13g2_buf_8
Xfanout2463 net2465 net2463 VPWR VGND sg13g2_buf_8
Xfanout2430 net2432 net2430 VPWR VGND sg13g2_buf_8
Xfanout2452 net2453 net2452 VPWR VGND sg13g2_buf_8
Xfanout2441 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2441 VPWR
+ VGND sg13g2_buf_8
XFILLER_78_762 VPWR VGND sg13g2_fill_1
XFILLER_66_913 VPWR VGND sg13g2_fill_1
Xfanout2496 net2497 net2496 VPWR VGND sg13g2_buf_8
Xfanout2485 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2485 VPWR VGND sg13g2_buf_8
Xfanout2474 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2474 VPWR
+ VGND sg13g2_buf_8
XFILLER_93_710 VPWR VGND sg13g2_fill_1
XFILLER_78_795 VPWR VGND sg13g2_fill_1
XFILLER_93_754 VPWR VGND sg13g2_decap_8
XFILLER_66_968 VPWR VGND sg13g2_fill_1
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_81_949 VPWR VGND sg13g2_decap_8
XFILLER_80_404 VPWR VGND sg13g2_fill_1
XFILLER_65_478 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2562 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_18_383 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q net3280 VGND VPWR i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[70\] clknet_leaf_75_clk sg13g2_dfrbpq_1
XFILLER_106_119 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2572 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2538 sg13g2_a21oi_1
XFILLER_1_909 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[357\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net828 net2447 net2272 VPWR VGND sg13g2_a22oi_1
XFILLER_103_837 VPWR VGND sg13g2_decap_8
XFILLER_102_336 VPWR VGND sg13g2_decap_8
XFILLER_29_38 VPWR VGND sg13g2_fill_1
XFILLER_84_710 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_xor2_1
Xdata_pdata\[4\]_sg13g2_mux2_1_A1 rsp_data_q\[4\] net698 net3051 data_pdata\[4\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_83_275 VPWR VGND sg13g2_decap_8
XFILLER_44_618 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2477 net2466 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_25_821 VPWR VGND sg13g2_fill_2
XFILLER_37_681 VPWR VGND sg13g2_decap_4
XFILLER_101_21 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_12_526 VPWR VGND sg13g2_decap_8
XFILLER_40_813 VPWR VGND sg13g2_decap_8
XFILLER_40_824 VPWR VGND sg13g2_fill_1
XFILLER_101_98 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[17\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.pc_d\[17\]
+ i_snitch.inst_addr_o\[17\] clknet_leaf_68_clk sg13g2_dfrbpq_2
XFILLER_4_725 VPWR VGND sg13g2_fill_1
XFILLER_106_631 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ net2523 VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.inst_addr_o\[25\] i_snitch.inst_addr_o\[26\] sg13g2_o21ai_1
XFILLER_105_196 VPWR VGND sg13g2_decap_8
XFILLER_79_559 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[4\] net1018 net2916 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_0_975 VPWR VGND sg13g2_decap_8
XFILLER_102_870 VPWR VGND sg13g2_decap_8
XFILLER_48_946 VPWR VGND sg13g2_decap_4
XFILLER_87_592 VPWR VGND sg13g2_decap_8
XFILLER_75_743 VPWR VGND sg13g2_fill_2
XFILLER_59_294 VPWR VGND sg13g2_decap_8
XFILLER_19_71 VPWR VGND sg13g2_fill_2
XFILLER_75_787 VPWR VGND sg13g2_fill_2
XFILLER_63_927 VPWR VGND sg13g2_decap_4
XFILLER_47_489 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[90\] clknet_leaf_111_clk sg13g2_dfrbpq_1
XFILLER_19_169 VPWR VGND sg13g2_decap_4
XFILLER_34_106 VPWR VGND sg13g2_fill_1
XFILLER_62_448 VPWR VGND sg13g2_fill_2
XFILLER_56_990 VPWR VGND sg13g2_fill_1
XFILLER_15_320 VPWR VGND sg13g2_fill_2
XFILLER_34_117 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q
+ net3245 VGND VPWR net1134 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_15_331 VPWR VGND sg13g2_fill_2
XFILLER_31_824 VPWR VGND sg13g2_fill_1
XFILLER_35_81 VPWR VGND sg13g2_fill_1
XFILLER_42_161 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y net2512
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[377\] clknet_leaf_114_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_xnor2_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nand2_1_B
+ target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[166\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2344 net1135 net2899 net2774 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\] net606 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xhold508 i_snitch.sb_q\[5\] VPWR VGND net540 sg13g2_dlygate4sd3_1
Xhold519 shift_reg_q\[26\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net551 sg13g2_dlygate4sd3_1
XFILLER_7_596 VPWR VGND sg13g2_fill_1
XFILLER_97_301 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2516 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2427 sg13g2_a21oi_1
XFILLER_98_857 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B_sg13g2_nand2_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B
+ net3076 net3075 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\] net2618 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xfanout2260 net2261 net2260 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ net2980 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net3008 i_snitch.sb_q\[1\] VPWR VGND sg13g2_a22oi_1
Xfanout2271 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2271 VPWR VGND sg13g2_buf_8
XFILLER_85_518 VPWR VGND sg13g2_fill_2
Xhold1208 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\] VPWR
+ VGND net1240 sg13g2_dlygate4sd3_1
Xfanout2293 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_Y
+ net2293 VPWR VGND sg13g2_buf_8
Xshift_reg_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2733 shift_reg_q\[18\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[14\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[14\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xfanout2282 net2283 net2282 VPWR VGND sg13g2_buf_8
Xhold1219 i_snitch.i_snitch_regfile.mem\[394\] VPWR VGND net1251 sg13g2_dlygate4sd3_1
XFILLER_38_434 VPWR VGND sg13g2_fill_1
XFILLER_65_253 VPWR VGND sg13g2_decap_8
XFILLER_25_106 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2706 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2613 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_30_890 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ net3078 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_1_706 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_89_846 VPWR VGND sg13g2_decap_8
XFILLER_88_301 VPWR VGND sg13g2_fill_1
XFILLER_0_216 VPWR VGND sg13g2_decap_8
XFILLER_102_133 VPWR VGND sg13g2_decap_8
XFILLER_88_345 VPWR VGND sg13g2_fill_1
XFILLER_0_249 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q
+ net3190 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[397\] clknet_leaf_85_clk sg13g2_dfrbpq_1
XFILLER_45_938 VPWR VGND sg13g2_fill_1
XFILLER_44_404 VPWR VGND sg13g2_decap_8
XFILLER_29_467 VPWR VGND sg13g2_decap_8
XFILLER_72_735 VPWR VGND sg13g2_fill_2
XFILLER_56_286 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[186\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2442 net2254 net2342 net1215 VPWR VGND sg13g2_a22oi_1
XFILLER_31_109 VPWR VGND sg13g2_fill_1
XFILLER_8_305 VPWR VGND sg13g2_fill_2
XFILLER_9_839 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a22oi_1_A1_Y
+ net2974 i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nand2b_1_A_N_Y net3006 i_snitch.i_snitch_regfile.mem\[34\]
+ VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2480 net2417 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y
+ net2498 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_450 VPWR VGND sg13g2_fill_1
XFILLER_97_21 VPWR VGND sg13g2_decap_8
XFILLER_97_98 VPWR VGND sg13g2_decap_4
XFILLER_79_356 VPWR VGND sg13g2_fill_1
XFILLER_0_772 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[35\]
+ net3006 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1_Y net2979 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[216\] clknet_leaf_57_clk sg13g2_dfrbpq_1
XFILLER_47_220 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_510 VPWR VGND sg13g2_decap_8
XFILLER_62_212 VPWR VGND sg13g2_decap_4
XFILLER_62_201 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1
+ VPWR VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_B2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2550 VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ VGND i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ net2715 sg13g2_o21ai_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]_sg13g2_nand2_1_B
+ i_req_register.data_o\[39\]_sg13g2_o21ai_1_Y_B1 net3173 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]
+ VPWR VGND sg13g2_nand2_1
Xstrb_reg_q\[5\]_sg13g2_a21oi_1_A1 VGND VPWR strb_reg_q\[5\] net3043 strb_reg_q\[5\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[4\]_sg13g2_a21oi_1_A1_B1 sg13g2_a21oi_1
XFILLER_30_153 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y net3007 sg13g2_o21ai_1
XFILLER_7_74 VPWR VGND sg13g2_fill_2
XFILLER_30_0 VPWR VGND sg13g2_fill_1
XFILLER_100_626 VPWR VGND sg13g2_decap_8
Xhold1005 i_snitch.i_snitch_regfile.mem\[92\] VPWR VGND net1037 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2844
+ sg13g2_a221oi_1
Xhold1027 i_snitch.i_snitch_regfile.mem\[119\] VPWR VGND net1059 sg13g2_dlygate4sd3_1
Xhold1016 i_snitch.i_snitch_regfile.mem\[192\] VPWR VGND net1048 sg13g2_dlygate4sd3_1
Xhold1049 i_snitch.i_snitch_regfile.mem\[303\] VPWR VGND net1081 sg13g2_dlygate4sd3_1
Xhold1038 i_snitch.i_snitch_regfile.mem\[339\] VPWR VGND net1070 sg13g2_dlygate4sd3_1
XFILLER_94_882 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_242 VPWR VGND sg13g2_decap_4
XFILLER_66_595 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_mux2_1_A0_X net3112 net2828 i_snitch.i_snitch_regfile.mem\[54\]
+ VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2_sg13g2_mux4_1_X
+ net3007 i_snitch.sb_q\[4\] i_snitch.sb_q\[5\] i_snitch.sb_q\[6\] i_snitch.sb_q\[7\]
+ net2980 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net1117 net2652 net2769 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2595 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_492 VPWR VGND sg13g2_decap_4
XFILLER_42_27 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_21_197 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B_sg13g2_nand3_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ net2933 net2941 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[236\] clknet_leaf_68_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_110_clk clknet_5_5__leaf_clk clknet_leaf_110_clk VPWR VGND sg13g2_buf_8
Xdata_pdata\[31\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2683 VPWR data_pdata\[31\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[31\]_sg13g2_nand2b_1_B_Y net3069 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1 net3000 i_snitch.i_snitch_regfile.mem\[410\]
+ i_snitch.i_snitch_regfile.mem\[442\] i_snitch.i_snitch_regfile.mem\[474\] i_snitch.i_snitch_regfile.mem\[506\]
+ net2976 i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] net601 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_104_921 VPWR VGND sg13g2_decap_8
XFILLER_89_610 VPWR VGND sg13g2_fill_1
Xhold861 i_snitch.inst_addr_o\[17\] VPWR VGND net893 sg13g2_dlygate4sd3_1
Xhold872 i_snitch.i_snitch_regfile.mem\[375\] VPWR VGND net904 sg13g2_dlygate4sd3_1
Xhold850 i_snitch.i_snitch_regfile.mem\[488\] VPWR VGND net882 sg13g2_dlygate4sd3_1
Xhold894 i_snitch.i_snitch_regfile.mem\[204\] VPWR VGND net926 sg13g2_dlygate4sd3_1
Xhold883 target_sel_q_sg13g2_nand2b_1_A_N_Y VPWR VGND net915 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_nand2_1_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_nand2_1_A_Y
+ net424 net2620 VPWR VGND sg13g2_nand2_1
XFILLER_104_998 VPWR VGND sg13g2_decap_8
XFILLER_103_486 VPWR VGND sg13g2_fill_1
XFILLER_88_175 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nor2_1_Y
+ net3076 net3075 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
XFILLER_76_337 VPWR VGND sg13g2_fill_1
XFILLER_76_326 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_85_871 VPWR VGND sg13g2_decap_8
XFILLER_29_264 VPWR VGND sg13g2_decap_8
XFILLER_83_34 VPWR VGND sg13g2_fill_1
XFILLER_17_437 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2604 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B
+ i_snitch.gpr_waddr\[7\]_sg13g2_nor2_1_A_Y data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_fill_1
XFILLER_13_654 VPWR VGND sg13g2_fill_2
XFILLER_34_1007 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.pc_d\[5\]
+ VGND net2301 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_8_135 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_101_clk clknet_5_19__leaf_clk clknet_leaf_101_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ sg13g2_o21ai_1
Xdata_pdata\[28\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[28\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[28\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
XFILLER_106_280 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y
+ VGND VPWR net2606 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_4_396 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\] net574 net2617
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net919 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2283
+ VPWR VGND sg13g2_a22oi_1
XFILLER_95_657 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_94_167 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net780 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2388 net3039 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
XFILLER_91_863 VPWR VGND sg13g2_decap_8
XFILLER_35_256 VPWR VGND sg13g2_decap_8
XFILLER_90_373 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[20\]_sg13g2_nor2_1_A net496 net2736 shift_reg_q\[20\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_63_598 VPWR VGND sg13g2_decap_4
XFILLER_23_429 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ net2716 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[75\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[75\]
+ net2846 i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q net3255 VGND VPWR i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[256\] clknet_leaf_106_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[423\]_sg13g2_o21ai_1_A1 net3091 VPWR i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[423\] net2810 sg13g2_o21ai_1
XFILLER_8_680 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1
+ net2600 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_mux2_1
XFILLER_104_217 VPWR VGND sg13g2_decap_8
XFILLER_99_930 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ net2708 sg13g2_or2_1
XFILLER_59_805 VPWR VGND sg13g2_fill_1
XFILLER_101_924 VPWR VGND sg13g2_decap_8
XFILLER_98_462 VPWR VGND sg13g2_fill_2
XFILLER_86_624 VPWR VGND sg13g2_decap_8
XFILLER_58_304 VPWR VGND sg13g2_fill_2
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.gpr_waddr\[7\]_sg13g2_nor2_1_A_Y
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2_X
+ VPWR VGND sg13g2_and2_1
XFILLER_100_456 VPWR VGND sg13g2_fill_1
XFILLER_67_871 VPWR VGND sg13g2_fill_1
XFILLER_66_370 VPWR VGND sg13g2_decap_8
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2419 sg13g2_a21oi_1
XFILLER_26_245 VPWR VGND sg13g2_decap_8
XFILLER_82_874 VPWR VGND sg13g2_decap_8
XFILLER_81_351 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C
+ net34 net48 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.wake_up_q\[2\]_sg13g2_nor4_1_D_Y_sg13g2_nand2_1_B i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B_Y
+ i_snitch.wake_up_q\[2\]_sg13g2_nor4_1_D_Y VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_23_952 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0_X
+ net3095 net2929 i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2641 i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_22_495 VPWR VGND sg13g2_fill_1
Xdata_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[4\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y data_pdata\[20\]_sg13g2_mux2_1_A0_X
+ net3153 sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net876 net2453 net2245 VPWR VGND sg13g2_a22oi_1
XFILLER_10_679 VPWR VGND sg13g2_fill_1
XFILLER_6_628 VPWR VGND sg13g2_fill_1
XFILLER_5_116 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
Xfanout2815 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X
+ net2815 VPWR VGND sg13g2_buf_8
XFILLER_89_440 VPWR VGND sg13g2_fill_1
Xhold680 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] VPWR
+ VGND net712 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2279
+ sg13g2_o21ai_1
Xfanout2837 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A
+ net2837 VPWR VGND sg13g2_buf_8
XFILLER_2_845 VPWR VGND sg13g2_decap_8
Xfanout2804 net2809 net2804 VPWR VGND sg13g2_buf_8
Xfanout2826 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_A2 net2826 VPWR
+ VGND sg13g2_buf_8
XFILLER_89_473 VPWR VGND sg13g2_fill_1
XFILLER_89_451 VPWR VGND sg13g2_fill_1
Xfanout2848 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y
+ net2848 VPWR VGND sg13g2_buf_8
Xhold691 i_snitch.i_snitch_regfile.mem\[337\] VPWR VGND net723 sg13g2_dlygate4sd3_1
Xfanout2859 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y
+ net2859 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ net2508 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_104_795 VPWR VGND sg13g2_decap_8
XFILLER_103_294 VPWR VGND sg13g2_decap_8
XFILLER_58_871 VPWR VGND sg13g2_decap_8
XFILLER_58_860 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q net3315 VGND VPWR i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[276\] clknet_leaf_66_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2459 net2855 i_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y net2309 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2 VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1
+ net2755 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_58_882 VPWR VGND sg13g2_fill_2
XFILLER_45_521 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1 net3015 i_snitch.i_snitch_regfile.mem\[414\]
+ i_snitch.i_snitch_regfile.mem\[446\] i_snitch.i_snitch_regfile.mem\[478\] i_snitch.i_snitch_regfile.mem\[510\]
+ net2985 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nand2_1_B_1
+ i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1_B1 net2972 net2958 VPWR VGND
+ sg13g2_nand2_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q
+ net3248 VGND VPWR net834 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2328
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A
+ net102 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_Y
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B VPWR
+ VGND sg13g2_or3_1
XFILLER_60_535 VPWR VGND sg13g2_decap_8
XFILLER_60_524 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ VGND net2604 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_14_974 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2591 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_43_92 VPWR VGND sg13g2_fill_1
XFILLER_9_411 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.sb_q\[11\] net2803 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_99_259 VPWR VGND sg13g2_fill_1
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_96_922 VPWR VGND sg13g2_decap_8
XFILLER_68_657 VPWR VGND sg13g2_decap_8
XFILLER_96_999 VPWR VGND sg13g2_decap_8
XFILLER_95_465 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_q\[12\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[12\] i_snitch.sb_q\[12\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_36_521 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_64_896 VPWR VGND sg13g2_decap_8
Xdata_pdata\[10\]_sg13g2_nand2b_1_B data_pdata\[10\]_sg13g2_nand2b_1_B_Y data_pdata\[10\]
+ net3157 VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y
+ net3080 i_req_arb.data_i\[44\] i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ net2720 sg13g2_a221oi_1
XFILLER_17_790 VPWR VGND sg13g2_fill_2
XFILLER_23_215 VPWR VGND sg13g2_fill_2
XFILLER_36_598 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2385
+ sg13g2_o21ai_1
XFILLER_104_1005 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B_sg13g2_nor2_1_Y
+ net2695 net2748 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_966 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and3_1_X
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_req_arb.data_i\[38\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ net2535 VPWR VGND sg13g2_and3_1
Xi_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q net3308 VGND VPWR i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[296\] clknet_leaf_70_clk sg13g2_dfrbpq_1
Xuo_out_sg13g2_buf_1_X_7 i_req_register.data_o\[41\] net24 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A
+ VPWR VGND sg13g2_nor3_1
XFILLER_87_944 VPWR VGND sg13g2_decap_8
XFILLER_86_410 VPWR VGND sg13g2_decap_8
XFILLER_59_624 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2731 shift_reg_q\[6\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[2\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_104_21 VPWR VGND sg13g2_decap_8
XFILLER_86_454 VPWR VGND sg13g2_fill_2
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_101_798 VPWR VGND sg13g2_decap_8
XFILLER_100_275 VPWR VGND sg13g2_decap_8
XFILLER_74_627 VPWR VGND sg13g2_decap_8
XFILLER_73_137 VPWR VGND sg13g2_fill_2
XFILLER_67_690 VPWR VGND sg13g2_fill_1
XFILLER_27_543 VPWR VGND sg13g2_fill_1
XFILLER_104_98 VPWR VGND sg13g2_decap_8
XFILLER_54_340 VPWR VGND sg13g2_decap_4
XFILLER_15_727 VPWR VGND sg13g2_decap_4
XFILLER_82_693 VPWR VGND sg13g2_fill_1
XFILLER_81_181 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nand2_1_A
+ i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A net1391 net3172
+ VPWR VGND sg13g2_nand2_2
XFILLER_27_598 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2415 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0 net3136 i_snitch.i_snitch_regfile.mem\[143\]
+ i_snitch.i_snitch_regfile.mem\[175\] i_snitch.i_snitch_regfile.mem\[207\] i_snitch.i_snitch_regfile.mem\[239\]
+ net3112 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xor2_1
XFILLER_22_281 VPWR VGND sg13g2_fill_1
XFILLER_7_948 VPWR VGND sg13g2_fill_1
XFILLER_6_458 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[115\] clknet_leaf_99_clk sg13g2_dfrbpq_1
Xfanout3313 net3329 net3313 VPWR VGND sg13g2_buf_8
Xfanout3302 net3306 net3302 VPWR VGND sg13g2_buf_8
Xfanout2601 net2602 net2601 VPWR VGND sg13g2_buf_1
Xfanout3324 net3325 net3324 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2259
+ sg13g2_o21ai_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2674 VPWR VGND sg13g2_nand2_1
XFILLER_2_642 VPWR VGND sg13g2_decap_8
Xfanout2612 net2615 net2612 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X
+ net51 net2848 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_Y
+ VPWR VGND sg13g2_nor4_1
Xfanout2634 net2636 net2634 VPWR VGND sg13g2_buf_8
Xfanout2623 net2624 net2623 VPWR VGND sg13g2_buf_8
Xfanout2645 net2646 net2645 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2921
+ sg13g2_a221oi_1
Xfanout2678 data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ net2678 VPWR VGND sg13g2_buf_8
Xdata_pdata\[30\]_sg13g2_nand2b_1_B data_pdata\[30\]_sg13g2_nand2b_1_B_Y data_pdata\[30\]
+ VPWR VGND net3162 sg13g2_nand2b_2
XFILLER_49_101 VPWR VGND sg13g2_fill_2
Xfanout2667 net2668 net2667 VPWR VGND sg13g2_buf_8
Xfanout2656 data_pdata\[28\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2656 VPWR
+ VGND sg13g2_buf_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2
+ net3073 net2926 VPWR VGND sg13g2_nand2_1
XFILLER_78_966 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ net2533 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y
+ net2482 VPWR VGND sg13g2_a22oi_1
Xfanout2689 data_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2689 VPWR VGND sg13g2_buf_8
XFILLER_93_958 VPWR VGND sg13g2_decap_8
XFILLER_77_476 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[14\]_sg13g2_dfrbpq_1_Q net3198 VGND VPWR net487 shift_reg_q\[14\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_64_137 VPWR VGND sg13g2_decap_4
XFILLER_18_521 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_45_362 VPWR VGND sg13g2_decap_4
XFILLER_61_844 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[483\]_sg13g2_o21ai_1_A1 net2962 VPWR i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[483\] net2801 sg13g2_o21ai_1
XFILLER_9_241 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0 net3014 i_snitch.i_snitch_regfile.mem\[262\]
+ i_snitch.i_snitch_regfile.mem\[294\] i_snitch.i_snitch_regfile.mem\[326\] i_snitch.i_snitch_regfile.mem\[358\]
+ net2986 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2252 net2387 net1176 VPWR VGND sg13g2_a22oi_1
XFILLER_86_1000 VPWR VGND sg13g2_decap_8
Xclkload22 clkload22/Y clknet_leaf_18_clk VPWR VGND sg13g2_inv_2
Xclkload11 clkload11/Y clknet_leaf_120_clk VPWR VGND sg13g2_inv_2
Xclkload33 VPWR clkload33/Y clknet_leaf_113_clk VGND sg13g2_inv_1
Xclkload44 clknet_leaf_76_clk clkload44/X VPWR VGND sg13g2_buf_8
Xclkload55 VPWR clkload55/Y clknet_leaf_54_clk VGND sg13g2_inv_1
Xclkload66 clkload66/Y clknet_leaf_56_clk VPWR VGND sg13g2_inv_2
XFILLER_6_970 VPWR VGND sg13g2_decap_8
XFILLER_102_507 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
XFILLER_69_922 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q_D VGND net310 net2322
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[82\]
+ i_snitch.i_snitch_regfile.mem\[114\] net3129 i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2694 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[272\] net3028 VPWR VGND sg13g2_nand2_1
XFILLER_84_947 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ net2586 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nand2b_1
XFILLER_83_446 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y VPWR
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ net2626 sg13g2_o21ai_1
XFILLER_37_841 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X net1378 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1
+ net2312 i_snitch.pc_d\[2\] VPWR VGND sg13g2_mux2_1
XFILLER_24_502 VPWR VGND sg13g2_fill_1
XFILLER_37_885 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_90_clk clknet_5_21__leaf_clk clknet_leaf_90_clk VPWR VGND sg13g2_buf_8
XFILLER_37_896 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q net3191 VGND VPWR i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[135\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_24_557 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_o21ai_1_A1 net2938 VPWR i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[302\] net2812 sg13g2_o21ai_1
XFILLER_51_387 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1226 net2495 net1233 VPWR VGND sg13g2_a22oi_1
Xclkload5 VPWR clkload5/Y clknet_leaf_0_clk VGND sg13g2_inv_1
XFILLER_20_730 VPWR VGND sg13g2_fill_1
XFILLER_20_752 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_Y i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_Y i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2860
+ net2897 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2968
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X
+ sg13g2_a221oi_1
XFILLER_105_301 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net457 net2395 VPWR VGND sg13g2_nand2_1
XFILLER_106_857 VPWR VGND sg13g2_decap_8
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
Xshift_reg_q\[2\]_sg13g2_a22oi_1_A1 uio_out_sg13g2_inv_1_Y_1_A shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 shift_reg_q\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_105_378 VPWR VGND sg13g2_decap_8
XFILLER_79_719 VPWR VGND sg13g2_fill_2
XFILLER_1_7 VPWR VGND sg13g2_decap_8
Xdata_pdata\[21\]_sg13g2_a21oi_1_A2 VGND VPWR net3155 data_pdata\[21\] data_pdata\[21\]_sg13g2_a21oi_1_A2_Y
+ net3150 sg13g2_a21oi_1
XFILLER_8_1011 VPWR VGND sg13g2_decap_8
XFILLER_87_741 VPWR VGND sg13g2_decap_8
XFILLER_101_562 VPWR VGND sg13g2_fill_2
XFILLER_86_273 VPWR VGND sg13g2_decap_8
XFILLER_74_413 VPWR VGND sg13g2_fill_1
XFILLER_19_318 VPWR VGND sg13g2_fill_2
Xdata_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[10\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[26\]_sg13g2_nand2b_1_B_Y net3150 data_pdata\[18\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[10\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
XFILLER_101_595 VPWR VGND sg13g2_fill_2
XFILLER_90_917 VPWR VGND sg13g2_decap_8
XFILLER_46_159 VPWR VGND sg13g2_fill_2
XFILLER_27_362 VPWR VGND sg13g2_decap_4
XFILLER_83_991 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[431\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net829 net2677 net2864 VPWR VGND sg13g2_a22oi_1
XFILLER_91_67 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_81_clk clknet_5_28__leaf_clk clknet_leaf_81_clk VPWR VGND sg13g2_buf_8
XFILLER_42_354 VPWR VGND sg13g2_decap_4
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.wake_up_q\[0\] clknet_leaf_36_clk sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_10_295 VPWR VGND sg13g2_decap_4
XFILLER_7_767 VPWR VGND sg13g2_decap_8
XFILLER_7_745 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2696 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2798
+ net2650 VPWR VGND sg13g2_nand2_1
Xfanout3121 net79 net3121 VPWR VGND sg13g2_buf_8
Xfanout3110 net3114 net3110 VPWR VGND sg13g2_buf_8
Xfanout3143 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1_X
+ net3143 VPWR VGND sg13g2_buf_8
Xfanout2420 net2421 net2420 VPWR VGND sg13g2_buf_2
Xfanout3154 net1403 net3154 VPWR VGND sg13g2_buf_8
XFILLER_3_962 VPWR VGND sg13g2_decap_8
Xfanout3165 net3167 net3165 VPWR VGND sg13g2_buf_8
Xfanout3132 net3132 net3140 VPWR VGND sg13g2_buf_16
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2554 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_97_549 VPWR VGND sg13g2_fill_2
XFILLER_97_527 VPWR VGND sg13g2_decap_8
Xfanout3176 net3176 net3183 VPWR VGND sg13g2_buf_16
Xfanout3198 net3200 net3198 VPWR VGND sg13g2_buf_8
Xfanout2442 net2444 net2442 VPWR VGND sg13g2_buf_8
Xfanout2431 net2432 net2431 VPWR VGND sg13g2_buf_8
Xfanout3187 net3188 net3187 VPWR VGND sg13g2_buf_8
Xfanout2453 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2453 VPWR
+ VGND sg13g2_buf_8
Xfanout2486 net2488 net2486 VPWR VGND sg13g2_buf_8
Xfanout2464 net2465 net2464 VPWR VGND sg13g2_buf_8
Xfanout2475 net2476 net2475 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ net2550 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
XFILLER_78_785 VPWR VGND sg13g2_fill_1
Xfanout2497 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_o21ai_1_A2_Y net2497 VPWR VGND
+ sg13g2_buf_8
Xi_snitch.gpr_waddr\[7\]_sg13g2_nor2b_1_A i_snitch.gpr_waddr\[7\] i_snitch.gpr_waddr\[6\]
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B VPWR
+ VGND sg13g2_nor2b_2
XFILLER_1_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q net3192 VGND VPWR i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[155\] clknet_leaf_119_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2461 VPWR VGND sg13g2_nand2_1
XFILLER_81_928 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_18_362 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2595 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_34_833 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_72_clk clknet_5_24__leaf_clk clknet_leaf_72_clk VPWR VGND sg13g2_buf_8
XFILLER_45_192 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A
+ net2546 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
XFILLER_61_674 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2934 i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2464
+ net2244 net2649 net2864 VPWR VGND sg13g2_a22oi_1
XFILLER_101_1008 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2879 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2
+ net2507 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_60_0 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ net2481 VPWR VGND sg13g2_a22oi_1
XFILLER_103_816 VPWR VGND sg13g2_decap_8
XFILLER_88_516 VPWR VGND sg13g2_decap_4
XFILLER_102_315 VPWR VGND sg13g2_decap_8
XFILLER_60_1014 VPWR VGND sg13g2_decap_8
XFILLER_96_582 VPWR VGND sg13g2_fill_1
XFILLER_69_774 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_57_958 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_X net3095 i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VPWR VGND
+ sg13g2_a22oi_1
XFILLER_28_148 VPWR VGND sg13g2_fill_2
XFILLER_71_416 VPWR VGND sg13g2_fill_2
XFILLER_71_427 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2881
+ net2654 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[195\]_sg13g2_nor3_1_A net1360 net2789 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xclkbuf_leaf_63_clk clknet_5_29__leaf_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_80_994 VPWR VGND sg13g2_decap_8
XFILLER_101_77 VPWR VGND sg13g2_decap_8
XFILLER_20_571 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[175\] clknet_leaf_81_clk sg13g2_dfrbpq_1
XFILLER_3_236 VPWR VGND sg13g2_decap_8
XFILLER_3_225 VPWR VGND sg13g2_decap_8
XFILLER_106_676 VPWR VGND sg13g2_decap_8
XFILLER_3_258 VPWR VGND sg13g2_fill_2
XFILLER_105_175 VPWR VGND sg13g2_decap_8
XFILLER_0_954 VPWR VGND sg13g2_decap_8
XFILLER_48_958 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[89\]
+ i_snitch.i_snitch_regfile.mem\[121\] net3119 i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_19_50 VPWR VGND sg13g2_decap_4
XFILLER_90_736 VPWR VGND sg13g2_fill_2
XFILLER_62_427 VPWR VGND sg13g2_decap_8
XFILLER_16_844 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1_1 VGND VPWR i_snitch.i_snitch_regfile.mem\[37\]
+ net3001 i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1_1_Y net2974 sg13g2_a21oi_1
XFILLER_27_170 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_54_clk clknet_5_26__leaf_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_15_387 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2783
+ net2674 VPWR VGND sg13g2_nand2_1
XFILLER_30_302 VPWR VGND sg13g2_fill_2
XFILLER_30_324 VPWR VGND sg13g2_decap_4
XFILLER_30_346 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[471\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2375 net716 net2647 net2743 VPWR VGND sg13g2_a22oi_1
Xhold509 shift_reg_q\[22\] VPWR VGND net541 sg13g2_dlygate4sd3_1
XFILLER_7_575 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0 net3007 i_snitch.i_snitch_regfile.mem\[388\]
+ i_snitch.i_snitch_regfile.mem\[420\] i_snitch.i_snitch_regfile.mem\[452\] i_snitch.i_snitch_regfile.mem\[484\]
+ net2980 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2815 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_98_836 VPWR VGND sg13g2_decap_8
Xfanout2261 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ net2261 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
Xfanout2250 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y
+ net2250 VPWR VGND sg13g2_buf_8
XFILLER_100_819 VPWR VGND sg13g2_decap_8
Xfanout2283 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y
+ net2283 VPWR VGND sg13g2_buf_8
Xfanout2272 net2273 net2272 VPWR VGND sg13g2_buf_8
Xhold1209 i_snitch.i_snitch_regfile.mem\[490\] VPWR VGND net1241 sg13g2_dlygate4sd3_1
Xfanout2294 net2295 net2294 VPWR VGND sg13g2_buf_8
XFILLER_66_733 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N_Y
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_53_405 VPWR VGND sg13g2_fill_2
Xdata_pdata\[16\]_sg13g2_mux2_1_A1 rsp_data_q\[16\] net809 net3050 data_pdata\[16\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_25_129 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[398\] net3028 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_45_clk clknet_5_15__leaf_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
XFILLER_53_449 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[195\] clknet_leaf_108_clk sg13g2_dfrbpq_1
XFILLER_61_482 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[501\] clknet_leaf_98_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[421\]_sg13g2_nor3_1_A net1328 net2860 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[43\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xoutput18 net18 uo_out[1] VPWR VGND sg13g2_buf_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X net1394 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1
+ net2313 i_snitch.pc_d\[20\] VPWR VGND sg13g2_mux2_1
XFILLER_102_112 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_97_880 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ net1170 VGND sg13g2_inv_1
XFILLER_102_189 VPWR VGND sg13g2_decap_8
XFILLER_99_1021 VPWR VGND sg13g2_decap_8
XFILLER_84_530 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[119\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net1059 net2648 net2871 VPWR VGND sg13g2_a22oi_1
XFILLER_56_210 VPWR VGND sg13g2_fill_1
XFILLER_57_777 VPWR VGND sg13g2_fill_2
XFILLER_57_766 VPWR VGND sg13g2_fill_2
XFILLER_56_232 VPWR VGND sg13g2_fill_1
XFILLER_84_585 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A
+ sg13g2_or2_1
Xclkbuf_leaf_36_clk clknet_5_10__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[491\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net1025 net2679 net2859 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_o21ai_1_A1 net3011 VPWR i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[39\] net2975 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_80_780 VPWR VGND sg13g2_fill_1
XFILLER_25_696 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2607 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[18\]_sg13g2_a22oi_1_A1 shift_reg_q\[18\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[18\] VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[20\]_sg13g2_mux2_1_A0 data_pdata\[20\] data_pdata\[28\] net3160 data_pdata\[20\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q
+ net3199 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
XFILLER_20_390 VPWR VGND sg13g2_fill_1
XFILLER_4_578 VPWR VGND sg13g2_fill_2
XFILLER_106_495 VPWR VGND sg13g2_decap_8
XFILLER_97_77 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[343\] VGND sg13g2_inv_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1 i_req_arb.gen_arbiter.rr_q VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y
+ VGND i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_A
+ sg13g2_o21ai_1
XFILLER_0_751 VPWR VGND sg13g2_decap_8
XFILLER_94_349 VPWR VGND sg13g2_fill_2
XFILLER_75_530 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 net2628 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_o21ai_1_A1 net2972 VPWR i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[382\] net2804 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3088 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ net2849 net3074 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ net2753 sg13g2_a221oi_1
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\] i_snitch.i_snitch_lsu.metadata_q\[0\] i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_Y
+ VPWR VGND data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y sg13g2_nand4_1
XFILLER_36_928 VPWR VGND sg13g2_decap_4
XFILLER_63_725 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[310\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2652 net2780 net2318 net1152 VPWR VGND sg13g2_a22oi_1
XFILLER_47_298 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_27_clk clknet_5_8__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_71_780 VPWR VGND sg13g2_fill_1
XFILLER_62_268 VPWR VGND sg13g2_decap_8
XFILLER_15_162 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[63\] clknet_leaf_71_clk sg13g2_dfrbpq_1
XFILLER_15_195 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2701 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2b_1
XFILLER_12_891 VPWR VGND sg13g2_decap_4
XFILLER_30_165 VPWR VGND sg13g2_fill_1
XFILLER_7_53 VPWR VGND sg13g2_decap_8
XFILLER_11_1019 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A_Y net2843 i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[311\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[311\]
+ net3019 i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_a21oi_1_A1_Y net2991 sg13g2_a21oi_1
XFILLER_7_361 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net1097 net2679 net2888 VPWR VGND sg13g2_a22oi_1
XFILLER_98_622 VPWR VGND sg13g2_decap_8
XFILLER_97_176 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold1006 i_snitch.i_snitch_regfile.mem\[91\] VPWR VGND net1038 sg13g2_dlygate4sd3_1
Xhold1017 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]
+ VPWR VGND net1049 sg13g2_dlygate4sd3_1
XFILLER_97_187 VPWR VGND sg13g2_decap_8
Xhold1028 i_snitch.i_snitch_regfile.mem\[116\] VPWR VGND net1060 sg13g2_dlygate4sd3_1
Xhold1039 i_snitch.i_snitch_regfile.mem\[59\] VPWR VGND net1071 sg13g2_dlygate4sd3_1
XFILLER_38_221 VPWR VGND sg13g2_fill_1
XFILLER_94_861 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A_sg13g2_and3_1_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ net3035 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ VPWR VGND sg13g2_and3_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.sb_q\[3\] i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_39_766 VPWR VGND sg13g2_fill_2
XFILLER_81_522 VPWR VGND sg13g2_fill_2
XFILLER_26_405 VPWR VGND sg13g2_fill_2
XFILLER_38_265 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B
+ net2631 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_81_533 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_18_clk clknet_5_12__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_26_449 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D_sg13g2_nor2b_1_Y
+ net3142 net3145 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D
+ VPWR VGND sg13g2_nor2b_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2531 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_and2_1_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_and2_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B
+ VGND VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ sg13g2_or2_1
Xdata_pdata\[4\]_sg13g2_dfrbpq_1_Q net3228 VGND VPWR net699 data_pdata\[4\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_21_165 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2711 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B_sg13g2_nor3_1_Y
+ net3 net1122 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nor3_1
Xshift_reg_q\[1\]_sg13g2_nor2_1_A net535 net2730 shift_reg_q\[1\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_104_900 VPWR VGND sg13g2_decap_8
XFILLER_101_7 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2843
+ sg13g2_a221oi_1
XFILLER_89_622 VPWR VGND sg13g2_fill_2
Xhold873 i_snitch.i_snitch_regfile.mem\[468\] VPWR VGND net905 sg13g2_dlygate4sd3_1
Xhold851 i_snitch.i_snitch_regfile.mem\[395\] VPWR VGND net883 sg13g2_dlygate4sd3_1
Xhold840 i_snitch.i_snitch_regfile.mem\[96\] VPWR VGND net872 sg13g2_dlygate4sd3_1
Xhold862 i_snitch.i_snitch_regfile.mem\[347\] VPWR VGND net894 sg13g2_dlygate4sd3_1
XFILLER_103_421 VPWR VGND sg13g2_decap_8
XFILLER_89_644 VPWR VGND sg13g2_fill_2
Xhold884 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net916 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_A1
+ net1166 VGND sg13g2_inv_1
Xhold895 data_pdata\[24\] VPWR VGND net927 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_nand2_1_B
+ i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_B1 net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[330\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2405 net997 net2473 net2282 VPWR VGND sg13g2_a22oi_1
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_104_977 VPWR VGND sg13g2_decap_8
XFILLER_88_143 VPWR VGND sg13g2_decap_4
XFILLER_77_817 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ net2511 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_103_498 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ VGND net2598 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_85_850 VPWR VGND sg13g2_decap_8
XFILLER_57_552 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2729 strb_reg_q\[4\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D strb_reg_q\[3\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[83\] clknet_leaf_100_clk sg13g2_dfrbpq_1
XFILLER_29_232 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2557 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_224 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2378
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2349 net924 net2645 net2887 VPWR VGND sg13g2_a22oi_1
XFILLER_9_604 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2722 i_snitch.inst_addr_o\[20\] sg13g2_a21oi_2
XFILLER_4_342 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_req_register.data_o\[40\]_sg13g2_mux2_1_X i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\] net3165 i_req_register.data_o\[40\]
+ VPWR VGND sg13g2_mux2_1
XFILLER_95_625 VPWR VGND sg13g2_decap_8
XFILLER_95_603 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2476 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_nor3_1_A_Y net2454 net2767 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_dfrbpq_1_Q_D
+ net2908 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_75_360 VPWR VGND sg13g2_fill_1
XFILLER_57_91 VPWR VGND sg13g2_decap_8
XFILLER_35_213 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2560 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_91_842 VPWR VGND sg13g2_decap_8
XFILLER_75_393 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xdata_pdata\[25\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[25\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[25\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
XFILLER_35_235 VPWR VGND sg13g2_decap_8
XFILLER_23_419 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2
+ net2942 net2953 VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[37\]_sg13g2_nor3_1_A net1340 net2765 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
XFILLER_31_430 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2405 net964 net2473 net2245 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X
+ VPWR VGND sg13g2_or4_1
Xclkbuf_leaf_7_clk clknet_5_2__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1
+ net2707 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2
+ net2614 VPWR VGND sg13g2_a22oi_1
XFILLER_101_903 VPWR VGND sg13g2_decap_8
XFILLER_99_986 VPWR VGND sg13g2_decap_8
XFILLER_98_452 VPWR VGND sg13g2_decap_4
XFILLER_59_839 VPWR VGND sg13g2_decap_8
XFILLER_86_658 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_X
+ net3093 net2931 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_96_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[179\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2442 net2270 net2342 net1259 VPWR VGND sg13g2_a22oi_1
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
XFILLER_39_596 VPWR VGND sg13g2_fill_1
XFILLER_93_190 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net831 net714 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_82_853 VPWR VGND sg13g2_decap_8
XFILLER_66_393 VPWR VGND sg13g2_fill_1
XFILLER_26_224 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[99\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[99\]
+ net2801 sg13g2_o21ai_1
XFILLER_42_706 VPWR VGND sg13g2_fill_2
XFILLER_54_599 VPWR VGND sg13g2_decap_4
XFILLER_53_49 VPWR VGND sg13g2_fill_2
XFILLER_53_38 VPWR VGND sg13g2_decap_8
Xdata_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[7\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y
+ data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y data_pdata\[31\]_sg13g2_a21oi_1_A2_Y
+ net3152 sg13g2_a21oi_2
XFILLER_10_625 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[19\] net745 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2415 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_2_824 VPWR VGND sg13g2_decap_8
Xi_req_register.data_o\[5\]_sg13g2_inv_1_A_Y_sg13g2_nor3_1_B state i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y
+ req_data_valid_sg13g2_o21ai_1_Y_B1 shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1 VPWR VGND
+ sg13g2_nor3_2
Xhold681 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net713 sg13g2_dlygate4sd3_1
Xhold670 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\] VPWR
+ VGND net702 sg13g2_dlygate4sd3_1
Xfanout2827 net2830 net2827 VPWR VGND sg13g2_buf_8
Xfanout2805 net2809 net2805 VPWR VGND sg13g2_buf_1
Xfanout2816 net2818 net2816 VPWR VGND sg13g2_buf_8
XFILLER_104_774 VPWR VGND sg13g2_decap_8
Xfanout2849 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X
+ net2849 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B
+ net2634 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xhold692 i_snitch.i_snitch_regfile.mem\[244\] VPWR VGND net724 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR net592 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[209\] clknet_leaf_82_clk sg13g2_dfrbpq_1
Xfanout2838 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A
+ net2838 VPWR VGND sg13g2_buf_8
XFILLER_103_273 VPWR VGND sg13g2_decap_8
XFILLER_89_496 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_92_606 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2574 VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VGND net2583 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_100_980 VPWR VGND sg13g2_decap_8
XFILLER_94_56 VPWR VGND sg13g2_decap_4
XFILLER_76_179 VPWR VGND sg13g2_fill_2
XFILLER_76_168 VPWR VGND sg13g2_fill_1
Xhold1370 i_snitch.gpr_waddr\[5\] VPWR VGND net1402 sg13g2_dlygate4sd3_1
XFILLER_94_89 VPWR VGND sg13g2_decap_8
XFILLER_45_555 VPWR VGND sg13g2_fill_1
XFILLER_72_374 VPWR VGND sg13g2_decap_8
XFILLER_45_577 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net986 net2470 net2272 VPWR VGND sg13g2_a22oi_1
XFILLER_32_205 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ VGND net2941 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2
+ sg13g2_o21ai_1
XFILLER_60_547 VPWR VGND sg13g2_fill_2
XFILLER_41_750 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y
+ VPWR VGND net3089 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1
+ net2634 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2496 net1387 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ net1378 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2417 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[371\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[371\]
+ net3116 i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_4_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[505\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2266 net2367 net1199 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[199\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net885 net2439 net2284 VPWR VGND sg13g2_a22oi_1
XFILLER_96_901 VPWR VGND sg13g2_decap_8
XFILLER_95_422 VPWR VGND sg13g2_fill_1
XFILLER_4_98 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_1 i_snitch.i_snitch_regfile.mem\[124\]
+ net2801 i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_1_Y VPWR VGND sg13g2_nor2_1
XFILLER_96_978 VPWR VGND sg13g2_decap_8
XFILLER_95_488 VPWR VGND sg13g2_decap_8
XFILLER_55_319 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[400\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_64_831 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net845 net2678 net2769 VPWR VGND sg13g2_a22oi_1
XFILLER_36_544 VPWR VGND sg13g2_fill_2
XFILLER_90_0 VPWR VGND sg13g2_decap_8
XFILLER_104_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A_sg13g2_nor4_1_Y net3
+ net553 net1122 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A VPWR VGND sg13g2_nor4_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2604 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[229\] clknet_leaf_4_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR net628 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
Xi_snitch.sb_q\[6\]_sg13g2_dfrbpq_1_Q net3250 VGND VPWR i_snitch.sb_d\[6\] i_snitch.sb_q\[6\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_105_527 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2340
+ sg13g2_o21ai_1
XFILLER_2_109 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y VPWR
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B
+ net2626 sg13g2_o21ai_1
XFILLER_87_923 VPWR VGND sg13g2_decap_8
XFILLER_101_722 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2358
+ sg13g2_o21ai_1
XFILLER_48_49 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2389 net1145 net2899 net3040 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR
+ VGND net2832 net2642 i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y net2955
+ i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y
+ sg13g2_a221oi_1
XFILLER_100_254 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and4_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net3036 net2927 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_and4_2
XFILLER_86_488 VPWR VGND sg13g2_decap_4
XFILLER_104_77 VPWR VGND sg13g2_decap_8
XFILLER_27_533 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2554 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2593 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2918
+ sg13g2_a221oi_1
XFILLER_11_956 VPWR VGND sg13g2_fill_1
Xfanout3303 net3306 net3303 VPWR VGND sg13g2_buf_8
Xfanout3314 net3316 net3314 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[420\] clknet_leaf_14_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xfanout2602 net2603 net2602 VPWR VGND sg13g2_buf_8
Xfanout3325 net3326 net3325 VPWR VGND sg13g2_buf_8
XFILLER_2_621 VPWR VGND sg13g2_decap_8
Xfanout2613 net2615 net2613 VPWR VGND sg13g2_buf_8
Xfanout2635 net2636 net2635 VPWR VGND sg13g2_buf_8
Xfanout2624 net2625 net2624 VPWR VGND sg13g2_buf_8
XFILLER_78_945 VPWR VGND sg13g2_decap_8
Xfanout2646 data_pdata\[31\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2646 VPWR
+ VGND sg13g2_buf_8
Xfanout2679 net2680 net2679 VPWR VGND sg13g2_buf_8
XFILLER_49_113 VPWR VGND sg13g2_fill_2
Xfanout2657 net2658 net2657 VPWR VGND sg13g2_buf_8
XFILLER_2_698 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_nand2_1_A_1 i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_nand2_1_A_1_Y
+ i_snitch.i_snitch_regfile.mem\[306\] net3016 VPWR VGND sg13g2_nand2_1
Xfanout2668 data_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2668 VPWR
+ VGND sg13g2_buf_8
XFILLER_93_937 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_and4_1_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B
+ VPWR VGND sg13g2_and4_1
XFILLER_65_617 VPWR VGND sg13g2_decap_4
XFILLER_92_436 VPWR VGND sg13g2_fill_2
XFILLER_46_831 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_57_190 VPWR VGND sg13g2_fill_1
XFILLER_45_385 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[249\] clknet_leaf_116_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ VGND net2707 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ sg13g2_o21ai_1
XFILLER_72_193 VPWR VGND sg13g2_decap_8
XFILLER_13_260 VPWR VGND sg13g2_fill_1
XFILLER_14_772 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] net653 net2624
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_13_282 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2745 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1
+ VGND VPWR net35 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ net112 net113 sg13g2_a21oi_2
Xclkload23 clkload23/Y clknet_leaf_23_clk VPWR VGND sg13g2_inv_2
XFILLER_9_297 VPWR VGND sg13g2_fill_1
Xclkload12 clkload12/Y clknet_leaf_110_clk VPWR VGND sg13g2_inv_2
Xclkload34 clknet_leaf_100_clk clkload34/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[100\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[100\]
+ net2803 sg13g2_o21ai_1
Xclkload67 clkload67/Y clknet_leaf_59_clk VPWR VGND sg13g2_inv_2
Xclkload56 clkload56/Y clknet_leaf_66_clk VPWR VGND sg13g2_inv_2
Xclkload45 clknet_leaf_77_clk clkload45/X VPWR VGND sg13g2_buf_8
XFILLER_5_481 VPWR VGND sg13g2_fill_1
XFILLER_5_470 VPWR VGND sg13g2_fill_2
XFILLER_48_2 VPWR VGND sg13g2_fill_1
XFILLER_96_720 VPWR VGND sg13g2_decap_4
XFILLER_68_411 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_96_764 VPWR VGND sg13g2_decap_8
XFILLER_84_926 VPWR VGND sg13g2_decap_8
XFILLER_68_466 VPWR VGND sg13g2_fill_1
XFILLER_95_285 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D
+ sg13g2_nand4_1
XFILLER_64_694 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2607 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ VGND net2718 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[440\] clknet_leaf_67_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2562 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[87\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net939 net2648 net2787 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_nor2_1_B
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nor2_1
Xclkload6 VPWR clkload6/Y clknet_leaf_5_clk VGND sg13g2_inv_1
Xrsp_state_q_sg13g2_dfrbpq_1_Q net3232 VGND VPWR rsp_state_d rsp_state_q clknet_leaf_36_clk
+ sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_106_836 VPWR VGND sg13g2_decap_8
XFILLER_105_357 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2886
+ net2669 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2558 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_101_541 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[269\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_101_585 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_75_937 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y
+ VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C
+ VGND i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B
+ net2576 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q
+ net3245 VGND VPWR net1090 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2792
+ net2693 VPWR VGND sg13g2_nand2_1
XFILLER_83_970 VPWR VGND sg13g2_decap_8
XFILLER_74_469 VPWR VGND sg13g2_fill_2
XFILLER_55_661 VPWR VGND sg13g2_fill_2
XFILLER_61_119 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2_1_A
+ net1391 net3164 req_data_valid_sg13g2_o21ai_1_Y_B1 VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2547 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xrsp_data_q\[21\]_sg13g2_dfrbpq_1_Q net3232 VGND VPWR rsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[21\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_10_252 VPWR VGND sg13g2_fill_1
XFILLER_10_285 VPWR VGND sg13g2_fill_1
Xfanout3111 net3114 net3111 VPWR VGND sg13g2_buf_8
Xfanout3122 net3125 net3122 VPWR VGND sg13g2_buf_8
Xfanout3100 net3101 net3100 VPWR VGND sg13g2_buf_8
Xfanout3144 net3146 net3144 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
Xfanout3133 net107 net3133 VPWR VGND sg13g2_buf_8
XFILLER_3_941 VPWR VGND sg13g2_decap_8
Xfanout3155 net3158 net3155 VPWR VGND sg13g2_buf_8
Xfanout2410 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y
+ net2410 VPWR VGND sg13g2_buf_8
Xfanout3177 net105 net3177 VPWR VGND sg13g2_buf_8
XFILLER_78_731 VPWR VGND sg13g2_fill_2
XFILLER_69_219 VPWR VGND sg13g2_decap_8
Xfanout2421 net2422 net2421 VPWR VGND sg13g2_buf_1
Xfanout2443 net2444 net2443 VPWR VGND sg13g2_buf_8
Xfanout3188 net3194 net3188 VPWR VGND sg13g2_buf_8
Xfanout3166 net3167 net3166 VPWR VGND sg13g2_buf_8
Xfanout2432 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2432 VPWR
+ VGND sg13g2_buf_8
Xfanout3199 net3200 net3199 VPWR VGND sg13g2_buf_8
Xfanout2487 net2488 net2487 VPWR VGND sg13g2_buf_1
Xfanout2454 net2455 net2454 VPWR VGND sg13g2_buf_8
Xfanout2465 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2465 VPWR
+ VGND sg13g2_buf_8
Xfanout2476 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2476 VPWR VGND sg13g2_buf_8
XFILLER_65_414 VPWR VGND sg13g2_fill_2
Xfanout2498 net2502 net2498 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2476 net2472 i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[460\] clknet_leaf_69_clk sg13g2_dfrbpq_1
XFILLER_81_907 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_18_330 VPWR VGND sg13g2_fill_2
XFILLER_33_300 VPWR VGND sg13g2_fill_2
XFILLER_73_491 VPWR VGND sg13g2_decap_8
XFILLER_21_517 VPWR VGND sg13g2_fill_1
XFILLER_14_591 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[289\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q
+ net3184 VGND VPWR net590 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
Xrsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2638 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1_X net2967 VPWR VGND sg13g2_a22oi_1
XFILLER_57_915 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[334\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2437
+ net2513 net2901 net2875 VPWR VGND sg13g2_a22oi_1
XFILLER_25_823 VPWR VGND sg13g2_fill_1
XFILLER_52_653 VPWR VGND sg13g2_decap_4
XFILLER_101_56 VPWR VGND sg13g2_decap_8
XFILLER_80_973 VPWR VGND sg13g2_decap_8
XFILLER_25_889 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[108\] clknet_leaf_71_clk sg13g2_dfrbpq_1
XFILLER_106_600 VPWR VGND sg13g2_fill_2
XFILLER_106_655 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[480\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_105_154 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A_Y net3012 sg13g2_o21ai_1
XFILLER_0_933 VPWR VGND sg13g2_decap_8
XFILLER_47_414 VPWR VGND sg13g2_fill_2
XFILLER_101_371 VPWR VGND sg13g2_decap_8
XFILLER_87_583 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X
+ net3076 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[154\]
+ i_snitch.i_snitch_regfile.mem\[186\] i_snitch.i_snitch_regfile.mem\[218\] i_snitch.i_snitch_regfile.mem\[250\]
+ net3098 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_75_767 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2543 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
XFILLER_76_1011 VPWR VGND sg13g2_decap_8
XFILLER_15_300 VPWR VGND sg13g2_decap_8
XFILLER_27_160 VPWR VGND sg13g2_decap_4
XFILLER_28_694 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_71_962 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2898 VPWR VGND sg13g2_nand2_1
XFILLER_42_130 VPWR VGND sg13g2_fill_2
XFILLER_70_472 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[270\]
+ net3028 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_a21oi_1_A1_Y net2988 sg13g2_a21oi_1
XFILLER_37_1017 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B
+ net109 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net1111 net2672 net3041 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[22\]_sg13g2_dfrbpq_1_Q net3204 VGND VPWR net799 data_pdata\[22\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_7_532 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2881
+ net2668 VPWR VGND sg13g2_nand2_1
XFILLER_98_815 VPWR VGND sg13g2_decap_8
XFILLER_83_1026 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2709 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xfanout2240 net2240 net68 VPWR VGND sg13g2_buf_16
Xfanout2251 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y
+ net2251 VPWR VGND sg13g2_buf_8
Xfanout2262 net2263 net2262 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_and2_1
XFILLER_78_550 VPWR VGND sg13g2_fill_1
Xfanout2295 net2298 net2295 VPWR VGND sg13g2_buf_8
Xfanout2284 net2285 net2284 VPWR VGND sg13g2_buf_8
Xfanout2273 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ net2273 VPWR VGND sg13g2_buf_8
XFILLER_39_948 VPWR VGND sg13g2_fill_1
XFILLER_81_748 VPWR VGND sg13g2_decap_8
XFILLER_81_737 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y VGND
+ VPWR net2615 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_62_962 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[128\] clknet_leaf_18_clk sg13g2_dfrbpq_1
Xshift_reg_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2731 shift_reg_q\[19\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[15\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[15\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_90_1008 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[93\]
+ i_snitch.i_snitch_regfile.mem\[125\] net3126 i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_A2
+ VGND VPWR net2584 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ net2579 sg13g2_a21oi_1
Xshift_reg_q\[27\]_sg13g2_dfrbpq_1_Q net3199 VGND VPWR net615 shift_reg_q\[27\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
Xoutput19 net19 uo_out[2] VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2777
+ net2898 VPWR VGND sg13g2_nand2_1
XFILLER_103_603 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2439 net2788 i_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2
+ net3034 net2927 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[326\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[326\] net2950 VPWR VGND sg13g2_nand2_1
XFILLER_102_168 VPWR VGND sg13g2_decap_8
XFILLER_69_572 VPWR VGND sg13g2_decap_4
XFILLER_99_1000 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0 net3133 i_snitch.i_snitch_regfile.mem\[392\]
+ i_snitch.i_snitch_regfile.mem\[424\] i_snitch.i_snitch_regfile.mem\[456\] i_snitch.i_snitch_regfile.mem\[488\]
+ net3113 i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_5_1026 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[290\]
+ net3002 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1_Y net2975 sg13g2_a21oi_1
XFILLER_29_414 VPWR VGND sg13g2_decap_8
XFILLER_84_597 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[424\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net816 net2644 net2863 VPWR VGND sg13g2_a22oi_1
XFILLER_38_981 VPWR VGND sg13g2_fill_1
XFILLER_72_59 VPWR VGND sg13g2_decap_8
XFILLER_52_450 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2
+ VGND i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_13_826 VPWR VGND sg13g2_decap_8
XFILLER_24_185 VPWR VGND sg13g2_decap_8
XFILLER_8_307 VPWR VGND sg13g2_fill_1
Xdata_pdata\[20\]_sg13g2_mux2_1_A1 net907 net925 net3050 data_pdata\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_380 VPWR VGND sg13g2_fill_2
XFILLER_106_441 VPWR VGND sg13g2_decap_8
XFILLER_97_56 VPWR VGND sg13g2_decap_8
XFILLER_79_336 VPWR VGND sg13g2_fill_1
XFILLER_79_325 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[148\] clknet_leaf_60_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2829
+ sg13g2_a221oi_1
XFILLER_0_730 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ net2429 VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2489 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ VPWR VGND sg13g2_and4_2
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[315\] net2810 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[445\] net3015 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[292\]_sg13g2_nor3_1_A net1320 net2778 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_94_328 VPWR VGND sg13g2_fill_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1
+ VPWR VGND sg13g2_and4_1
XFILLER_47_255 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2768
+ net2676 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ net2580 sg13g2_or2_1
XFILLER_29_981 VPWR VGND sg13g2_fill_2
XFILLER_35_406 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ sg13g2_o21ai_1
Xshift_reg_q\[15\]_sg13g2_nor2_1_A net461 net2732 shift_reg_q\[15\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_675 VPWR VGND sg13g2_fill_2
XFILLER_94_7 VPWR VGND sg13g2_decap_8
XFILLER_43_472 VPWR VGND sg13g2_fill_2
XFILLER_70_291 VPWR VGND sg13g2_fill_2
XFILLER_30_133 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2892
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_50_1025 VPWR VGND sg13g2_decap_4
XFILLER_30_177 VPWR VGND sg13g2_fill_2
XFILLER_8_852 VPWR VGND sg13g2_fill_2
XFILLER_7_32 VPWR VGND sg13g2_decap_8
XFILLER_30_199 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[444\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2464 net2246 net2381 net1202 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2778 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2910 net678 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D net2320
+ sg13g2_a221oi_1
XFILLER_98_678 VPWR VGND sg13g2_decap_8
XFILLER_85_317 VPWR VGND sg13g2_fill_2
Xhold1018 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1050 sg13g2_dlygate4sd3_1
Xhold1029 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]
+ VPWR VGND net1061 sg13g2_dlygate4sd3_1
Xhold1007 i_snitch.i_snitch_regfile.mem\[209\] VPWR VGND net1039 sg13g2_dlygate4sd3_1
XFILLER_94_840 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
XFILLER_27_907 VPWR VGND sg13g2_decap_4
XFILLER_39_756 VPWR VGND sg13g2_decap_4
XFILLER_54_759 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2845
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] net3179 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_50_943 VPWR VGND sg13g2_fill_2
Xdata_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2714 data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y net3070 sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xdata_pvalid_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y net1408 net2488 data_pvalid_sg13g2_nor2_1_A_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_a21oi_1_A1_Y net2642 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y
+ net2955 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[168\] clknet_leaf_73_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net2695 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1
+ sg13g2_a21oi_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2630 net2760 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_a22oi_1
Xhold830 i_snitch.i_snitch_regfile.mem\[472\] VPWR VGND net862 sg13g2_dlygate4sd3_1
Xhold841 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] VPWR
+ VGND net873 sg13g2_dlygate4sd3_1
Xhold863 i_snitch.i_snitch_regfile.mem\[367\] VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold852 i_snitch.i_snitch_regfile.mem\[285\] VPWR VGND net884 sg13g2_dlygate4sd3_1
XFILLER_104_956 VPWR VGND sg13g2_decap_8
XFILLER_89_656 VPWR VGND sg13g2_fill_2
Xhold885 i_snitch.i_snitch_regfile.mem\[287\] VPWR VGND net917 sg13g2_dlygate4sd3_1
Xhold896 data_pdata\[24\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net928 sg13g2_dlygate4sd3_1
Xhold874 i_snitch.i_snitch_regfile.mem\[175\] VPWR VGND net906 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2749 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_89_689 VPWR VGND sg13g2_fill_2
XFILLER_89_678 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2479 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y
+ net2530 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2
+ net2546 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2378
+ sg13g2_o21ai_1
XFILLER_45_759 VPWR VGND sg13g2_decap_4
XFILLER_52_280 VPWR VGND sg13g2_decap_4
XFILLER_25_483 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2597 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_40_442 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[464\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net983 net2461 net2262 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B_Y i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2919
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C i_snitch.inst_addr_o\[25\]
+ net2305 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_10_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_79_188 VPWR VGND sg13g2_fill_1
XFILLER_48_520 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y net3020 sg13g2_o21ai_1
XFILLER_48_531 VPWR VGND sg13g2_decap_8
XFILLER_63_501 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2962
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A net2963
+ net2958 VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0 net3135 i_snitch.i_snitch_regfile.mem\[399\]
+ i_snitch.i_snitch_regfile.mem\[431\] i_snitch.i_snitch_regfile.mem\[463\] i_snitch.i_snitch_regfile.mem\[495\]
+ net3112 i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_17_940 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X
+ net2684 net2746 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_mux2_1
XFILLER_91_898 VPWR VGND sg13g2_decap_8
XFILLER_90_364 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[188\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2627 net2851 net3082
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_965 VPWR VGND sg13g2_decap_8
XFILLER_89_1021 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_dfrbpq_1_Q net3224 VGND VPWR i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[36\] clknet_leaf_107_clk sg13g2_dfrbpq_1
Xdata_pdata\[27\]_sg13g2_mux2_1_A1 rsp_data_q\[27\] net941 net3049 data_pdata\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_99_965 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y
+ net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\] VPWR
+ VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_101_959 VPWR VGND sg13g2_decap_8
XFILLER_100_425 VPWR VGND sg13g2_fill_2
XFILLER_98_497 VPWR VGND sg13g2_fill_2
XFILLER_98_486 VPWR VGND sg13g2_decap_4
XFILLER_58_339 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y
+ net2746 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_82_810 VPWR VGND sg13g2_fill_1
XFILLER_67_884 VPWR VGND sg13g2_fill_2
Xstrb_reg_q\[6\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ strb_reg_q\[6\] clknet_leaf_122_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[14\] net1089 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_81_386 VPWR VGND sg13g2_decap_8
XFILLER_34_280 VPWR VGND sg13g2_fill_2
XFILLER_50_795 VPWR VGND sg13g2_fill_2
XFILLER_23_998 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q
+ net3231 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_10_637 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_inv_1_A
+ net860 i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_A2 VPWR VGND sg13g2_inv_4
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net88 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xrebuffer278 net310 net2257 VPWR VGND sg13g2_buf_16
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2501 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[485\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[485\]
+ net3117 i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_2_803 VPWR VGND sg13g2_decap_8
Xfanout2806 net2807 net2806 VPWR VGND sg13g2_buf_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
Xfanout2828 net2829 net2828 VPWR VGND sg13g2_buf_8
Xhold660 i_snitch.i_snitch_lsu.metadata_q\[9\] VPWR VGND net692 sg13g2_dlygate4sd3_1
Xhold671 i_snitch.i_snitch_regfile.mem\[346\] VPWR VGND net703 sg13g2_dlygate4sd3_1
Xfanout2817 net2818 net2817 VPWR VGND sg13g2_buf_2
XFILLER_103_252 VPWR VGND sg13g2_decap_8
Xhold682 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\] VPWR
+ VGND net714 sg13g2_dlygate4sd3_1
Xfanout2839 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A
+ net2839 VPWR VGND sg13g2_buf_8
Xhold693 data_pdata\[13\] VPWR VGND net725 sg13g2_dlygate4sd3_1
Xdata_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y data_pdata\[21\]_sg13g2_mux2_1_A0_X
+ net3151 sg13g2_a21oi_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_2
Xi_snitch.i_snitch_regfile.mem\[375\]_sg13g2_o21ai_1_A1 net2972 VPWR i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[375\] net2808 sg13g2_o21ai_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_94_35 VPWR VGND sg13g2_decap_8
XFILLER_76_136 VPWR VGND sg13g2_fill_2
Xhold1360 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A VPWR
+ VGND net1392 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_a22oi_1_A1_Y
+ net2677 net2781 net2319 net1081 VPWR VGND sg13g2_a22oi_1
Xhold1371 i_snitch.i_snitch_lsu.metadata_q\[3\] VPWR VGND net1403 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q_D VGND net2315 net2299
+ sg13g2_o21ai_1
XFILLER_17_247 VPWR VGND sg13g2_fill_1
XFILLER_33_718 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[56\] clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_14_921 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2419 sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X
+ net3072 i_snitch.sb_q\[4\] i_snitch.sb_q\[5\] i_snitch.sb_q\[6\] i_snitch.sb_q\[7\]
+ net3071 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[164\]_sg13g2_nor3_1_A net1290 net2776 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_40_283 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2328
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[304\]
+ net3016 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_a21oi_1_A1_Y net2987 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2476 i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2448 net2867 i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q_D net2908
+ sg13g2_a221oi_1
XFILLER_57_7 VPWR VGND sg13g2_decap_4
XFILLER_5_663 VPWR VGND sg13g2_fill_1
XFILLER_4_140 VPWR VGND sg13g2_decap_8
XFILLER_99_239 VPWR VGND sg13g2_fill_2
XFILLER_68_604 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
Xdata_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[1\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y
+ data_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y data_pdata\[25\]_sg13g2_a21oi_1_A2_Y
+ net3149 sg13g2_a21oi_2
XFILLER_96_957 VPWR VGND sg13g2_decap_8
XFILLER_83_629 VPWR VGND sg13g2_decap_8
XFILLER_64_821 VPWR VGND sg13g2_fill_1
XFILLER_49_895 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3092 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2377
+ sg13g2_o21ai_1
XFILLER_51_526 VPWR VGND sg13g2_decap_4
XFILLER_17_770 VPWR VGND sg13g2_decap_8
XFILLER_23_217 VPWR VGND sg13g2_fill_1
XFILLER_36_589 VPWR VGND sg13g2_fill_1
XFILLER_90_194 VPWR VGND sg13g2_decap_4
XFILLER_83_0 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_o21ai_1_A1 net3097 VPWR i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[395\] i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2515 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2427 sg13g2_a21oi_1
XFILLER_99_762 VPWR VGND sg13g2_decap_4
XFILLER_87_902 VPWR VGND sg13g2_decap_8
Xi_req_arb.data_i\[41\]_sg13g2_a21oi_1_B1 VGND VPWR net3086 net2536 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A
+ i_req_arb.data_i\[41\] sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2533 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ net2482 VPWR VGND sg13g2_a22oi_1
XFILLER_63_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y VGND
+ VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net54 net2611 sg13g2_a21oi_2
XFILLER_59_626 VPWR VGND sg13g2_fill_1
XFILLER_100_233 VPWR VGND sg13g2_decap_8
XFILLER_87_979 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q net3310 VGND VPWR i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[76\] clknet_leaf_69_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2347
+ sg13g2_o21ai_1
XFILLER_104_56 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_nand2b_1_A_N_Y
+ net3027 i_snitch.i_snitch_regfile.mem\[85\] VPWR VGND sg13g2_nand2b_1
XFILLER_27_523 VPWR VGND sg13g2_fill_1
XFILLER_70_813 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
Xshift_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2732 shift_reg_q\[7\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[3\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_42_515 VPWR VGND sg13g2_fill_1
XFILLER_42_526 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2364
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2595 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ net2587 sg13g2_a21oi_1
XFILLER_22_272 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A i_snitch.pc_d\[22\]_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[22\] VPWR VGND sg13g2_and2_1
XFILLER_6_405 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor3_1_C
+ net2567 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2392
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y
+ net3146 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1
+ VPWR VGND sg13g2_nand2_1
Xfanout3304 net3306 net3304 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]
+ net118 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
Xfanout3326 net3329 net3326 VPWR VGND sg13g2_buf_8
Xfanout3315 net3316 net3315 VPWR VGND sg13g2_buf_1
XFILLER_2_600 VPWR VGND sg13g2_decap_8
Xfanout2603 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y
+ net2603 VPWR VGND sg13g2_buf_8
Xfanout2614 net2615 net2614 VPWR VGND sg13g2_buf_1
Xfanout2636 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y
+ net2636 VPWR VGND sg13g2_buf_8
Xfanout2625 target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B_Y net2625
+ VPWR VGND sg13g2_buf_8
Xhold490 shift_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net522 sg13g2_dlygate4sd3_1
XFILLER_77_412 VPWR VGND sg13g2_fill_1
Xfanout2647 data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2647 VPWR
+ VGND sg13g2_buf_8
Xfanout2669 net2670 net2669 VPWR VGND sg13g2_buf_8
XFILLER_2_677 VPWR VGND sg13g2_decap_8
Xfanout2658 data_pdata\[27\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y net2658 VPWR
+ VGND sg13g2_buf_8
XFILLER_93_916 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2248
+ sg13g2_o21ai_1
XFILLER_38_50 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[325\] VGND sg13g2_inv_1
XFILLER_73_651 VPWR VGND sg13g2_fill_2
XFILLER_61_813 VPWR VGND sg13g2_fill_1
XFILLER_61_802 VPWR VGND sg13g2_fill_1
Xhold1190 i_snitch.i_snitch_regfile.mem\[507\] VPWR VGND net1222 sg13g2_dlygate4sd3_1
XFILLER_14_762 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[343\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2403 net891 net2647 net2796 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2573 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ net2538 sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A
+ net114 net3075 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q net3257 VGND VPWR i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[96\] clknet_leaf_49_clk sg13g2_dfrbpq_1
Xclkload24 VPWR clkload24/Y clknet_leaf_17_clk VGND sg13g2_inv_1
Xclkload35 clknet_leaf_104_clk clkload35/Y VPWR VGND sg13g2_inv_4
Xclkload13 clknet_leaf_14_clk clkload13/X VPWR VGND sg13g2_buf_8
Xclkload57 VPWR clkload57/Y clknet_leaf_68_clk VGND sg13g2_inv_1
XFILLER_55_4 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2531 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X
+ net2480 VPWR VGND sg13g2_a22oi_1
Xclkload46 VPWR clkload46/Y clknet_leaf_78_clk VGND sg13g2_inv_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 net2629
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2b_1
XFILLER_69_913 VPWR VGND sg13g2_fill_1
XFILLER_96_710 VPWR VGND sg13g2_decap_4
XFILLER_96_743 VPWR VGND sg13g2_decap_8
XFILLER_95_242 VPWR VGND sg13g2_decap_8
XFILLER_84_905 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_96_776 VPWR VGND sg13g2_fill_2
XFILLER_49_670 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2790 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2
+ net2504 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
Xrsp_data_q\[2\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR rsp_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[2\] clknet_leaf_38_clk sg13g2_dfrbpq_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2596 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_93_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_20_721 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2790
+ i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xclkload7 clkload7/Y clknet_leaf_10_clk VPWR VGND sg13g2_inv_2
XFILLER_106_815 VPWR VGND sg13g2_decap_8
XFILLER_105_336 VPWR VGND sg13g2_decap_8
XFILLER_59_27 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q
+ net3195 VGND VPWR net631 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_87_710 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] net639 net2624
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2
+ net3072 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net3071 i_snitch.sb_q\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_101_520 VPWR VGND sg13g2_fill_1
XFILLER_86_231 VPWR VGND sg13g2_fill_2
XFILLER_59_456 VPWR VGND sg13g2_decap_4
XFILLER_101_564 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ net63 net2761 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[363\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net848 net2680 net2882 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1
+ VGND VPWR net2569 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ net90 sg13g2_a21oi_1
XFILLER_91_14 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1_sg13g2_nor3_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1
+ VPWR VGND sg13g2_nor3_1
XFILLER_15_504 VPWR VGND sg13g2_fill_2
XFILLER_42_301 VPWR VGND sg13g2_fill_2
XFILLER_42_334 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q net3204 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[2\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_30_518 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.sb_q\[15\] net3122 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2941 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2511 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[364\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[364\]
+ net3134 i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
Xfanout3112 net3114 net3112 VPWR VGND sg13g2_buf_8
XFILLER_3_920 VPWR VGND sg13g2_decap_8
Xfanout3101 net3102 net3101 VPWR VGND sg13g2_buf_8
Xfanout3145 net3146 net3145 VPWR VGND sg13g2_buf_8
Xfanout3134 net3140 net3134 VPWR VGND sg13g2_buf_8
Xfanout3123 net3125 net3123 VPWR VGND sg13g2_buf_8
Xfanout2400 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2400 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_1 i_snitch.i_snitch_regfile.mem\[117\]
+ net2802 i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_1_Y VPWR VGND sg13g2_nor2_1
Xfanout3156 net3157 net3156 VPWR VGND sg13g2_buf_1
Xfanout2411 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y
+ net2411 VPWR VGND sg13g2_buf_8
XFILLER_97_518 VPWR VGND sg13g2_decap_4
Xfanout3178 net3182 net3178 VPWR VGND sg13g2_buf_8
XFILLER_78_710 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\] data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y
+ VPWR VGND sg13g2_nand2_1
Xfanout2422 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2422 VPWR VGND sg13g2_buf_8
Xfanout2444 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2444 VPWR
+ VGND sg13g2_buf_8
XFILLER_3_997 VPWR VGND sg13g2_decap_8
Xfanout3167 net3173 net3167 VPWR VGND sg13g2_buf_8
Xfanout3189 net3193 net3189 VPWR VGND sg13g2_buf_8
Xfanout2433 net2435 net2433 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_1 i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_1_Y
+ net2994 i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_nand2b_1_A_N_Y net3022 i_snitch.i_snitch_regfile.mem\[55\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_2_496 VPWR VGND sg13g2_fill_2
Xfanout2455 net2456 net2455 VPWR VGND sg13g2_buf_8
Xfanout2477 net2478 net2477 VPWR VGND sg13g2_buf_8
Xfanout2466 net2468 net2466 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]
+ net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xfanout2488 i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y net2488 VPWR
+ VGND sg13g2_buf_8
Xfanout2499 net2502 net2499 VPWR VGND sg13g2_buf_8
XFILLER_38_607 VPWR VGND sg13g2_decap_4
XFILLER_93_746 VPWR VGND sg13g2_fill_2
XFILLER_1_56 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net110
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2704 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2b_1
XFILLER_92_278 VPWR VGND sg13g2_fill_2
XFILLER_73_481 VPWR VGND sg13g2_fill_1
XFILLER_45_150 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_dfrbpq_1_Q
+ net3199 VGND VPWR net659 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2542 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
XFILLER_88_529 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ net2526 VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.inst_addr_o\[21\] i_snitch.inst_addr_o\[22\] sg13g2_o21ai_1
XFILLER_69_710 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[383\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[383\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2394 net802 net2645 net2880 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1
+ net745 net564 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_84_735 VPWR VGND sg13g2_decap_8
XFILLER_56_437 VPWR VGND sg13g2_decap_4
XFILLER_83_234 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ net2581 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_nand2b_1
XFILLER_71_418 VPWR VGND sg13g2_fill_1
XFILLER_80_952 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A
+ sg13g2_o21ai_1
XFILLER_52_632 VPWR VGND sg13g2_decap_8
XFILLER_101_35 VPWR VGND sg13g2_decap_8
XFILLER_52_665 VPWR VGND sg13g2_decap_4
XFILLER_24_389 VPWR VGND sg13g2_decap_8
XFILLER_40_838 VPWR VGND sg13g2_fill_2
XFILLER_20_551 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[274\] net2814 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q net3270 VGND VPWR i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[413\] clknet_leaf_95_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]
+ net3167 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_105_133 VPWR VGND sg13g2_decap_8
XFILLER_10_54 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[202\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net913 net2440 net2282 VPWR VGND sg13g2_a22oi_1
XFILLER_10_87 VPWR VGND sg13g2_fill_2
XFILLER_0_912 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[101\]
+ net2947 i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2
+ net2505 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_86_47 VPWR VGND sg13g2_decap_8
XFILLER_86_36 VPWR VGND sg13g2_fill_2
XFILLER_101_350 VPWR VGND sg13g2_decap_8
XFILLER_75_713 VPWR VGND sg13g2_decap_8
XFILLER_47_404 VPWR VGND sg13g2_decap_4
XFILLER_0_989 VPWR VGND sg13g2_decap_8
XFILLER_102_884 VPWR VGND sg13g2_decap_8
XFILLER_75_724 VPWR VGND sg13g2_fill_2
XFILLER_19_41 VPWR VGND sg13g2_decap_4
XFILLER_74_256 VPWR VGND sg13g2_decap_4
XFILLER_74_245 VPWR VGND sg13g2_fill_1
XFILLER_56_960 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[83\] net2977 VPWR VGND sg13g2_nand2_1
XFILLER_90_738 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1_sg13g2_and4_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net3035 net3073 net2926 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1
+ VPWR VGND sg13g2_and4_1
XFILLER_55_492 VPWR VGND sg13g2_fill_1
XFILLER_27_172 VPWR VGND sg13g2_fill_1
XFILLER_70_462 VPWR VGND sg13g2_fill_1
XFILLER_70_451 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2934 i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
XFILLER_30_304 VPWR VGND sg13g2_fill_1
XFILLER_35_95 VPWR VGND sg13g2_fill_1
XFILLER_42_197 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2638 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_83_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_772 VPWR VGND sg13g2_decap_8
XFILLER_97_359 VPWR VGND sg13g2_decap_4
Xfanout2241 i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C_Y
+ net2241 VPWR VGND sg13g2_buf_8
Xshift_reg_q\[4\]_sg13g2_dfrbpq_1_Q net3227 VGND VPWR net466 shift_reg_q\[4\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
Xfanout2252 net2253 net2252 VPWR VGND sg13g2_buf_8
XFILLER_3_783 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B net2628
+ VPWR VGND sg13g2_nand2_1
Xfanout2285 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y
+ net2285 VPWR VGND sg13g2_buf_8
Xfanout2263 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y
+ net2263 VPWR VGND sg13g2_buf_8
Xfanout2274 net2275 net2274 VPWR VGND sg13g2_buf_8
Xfanout2296 net2297 net2296 VPWR VGND sg13g2_buf_8
XFILLER_93_554 VPWR VGND sg13g2_fill_1
XFILLER_66_768 VPWR VGND sg13g2_decap_8
XFILLER_65_234 VPWR VGND sg13g2_decap_8
XFILLER_54_919 VPWR VGND sg13g2_decap_4
XFILLER_47_960 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2885
+ net2673 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[294\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[294\] net2812 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[433\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_22_849 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[222\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net972 net2440 net2244 VPWR VGND sg13g2_a22oi_1
XFILLER_21_348 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_122_clk clknet_5_0__leaf_clk clknet_leaf_122_clk VPWR VGND sg13g2_buf_8
XFILLER_30_860 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2779
+ net2668 VPWR VGND sg13g2_nand2_1
XFILLER_102_147 VPWR VGND sg13g2_decap_8
XFILLER_5_1005 VPWR VGND sg13g2_decap_8
XFILLER_29_404 VPWR VGND sg13g2_fill_1
XFILLER_57_779 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.inst_addr_o\[13\] net2528 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ net2551 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2439 net2788 i_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
XFILLER_80_771 VPWR VGND sg13g2_fill_1
XFILLER_53_985 VPWR VGND sg13g2_fill_2
XFILLER_24_153 VPWR VGND sg13g2_decap_4
XFILLER_12_315 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[14\]_sg13g2_dfrbpq_1_Q net3241 VGND VPWR rsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[14\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A_Y
+ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_113_clk clknet_5_16__leaf_clk clknet_leaf_113_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[79\] VGND sg13g2_inv_1
XFILLER_106_420 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2774
+ net2675 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A
+ sg13g2_a21oi_1
XFILLER_97_35 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2873
+ net2897 VPWR VGND sg13g2_nand2_1
XFILLER_88_882 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_0_786 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[453\] clknet_leaf_110_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y net2512
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_63_727 VPWR VGND sg13g2_fill_1
XFILLER_63_716 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[242\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net1012 net2438 net2272 VPWR VGND sg13g2_a22oi_1
XFILLER_62_226 VPWR VGND sg13g2_decap_8
XFILLER_16_632 VPWR VGND sg13g2_fill_1
XFILLER_90_568 VPWR VGND sg13g2_decap_4
XFILLER_43_440 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1
+ VGND sg13g2_inv_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[330\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[330\] net2950 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VGND net2566 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C
+ net3077 net3079 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
XFILLER_7_11 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_104_clk clknet_5_18__leaf_clk clknet_leaf_104_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0 net3135 i_snitch.i_snitch_regfile.mem\[401\]
+ i_snitch.i_snitch_regfile.mem\[433\] i_snitch.i_snitch_regfile.mem\[465\] i_snitch.i_snitch_regfile.mem\[497\]
+ net3112 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y
+ net2565 net2548 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C
+ VPWR VGND sg13g2_nor2_1
Xshift_reg_q\[9\]_sg13g2_nor2_1_A net538 net2728 shift_reg_q\[9\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_o21ai_1_A1 net3107 VPWR i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[449\] net3128 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[127\]
+ net2802 i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q
+ net3238 VGND VPWR net1066 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_98_602 VPWR VGND sg13g2_fill_2
XFILLER_98_657 VPWR VGND sg13g2_fill_2
XFILLER_97_134 VPWR VGND sg13g2_decap_4
Xhold1019 rsp_data_q\[28\] VPWR VGND net1051 sg13g2_dlygate4sd3_1
XFILLER_79_893 VPWR VGND sg13g2_decap_8
Xhold1008 i_snitch.i_snitch_regfile.mem\[62\] VPWR VGND net1040 sg13g2_dlygate4sd3_1
XFILLER_38_212 VPWR VGND sg13g2_decap_4
XFILLER_66_532 VPWR VGND sg13g2_decap_8
XFILLER_94_896 VPWR VGND sg13g2_decap_8
XFILLER_38_267 VPWR VGND sg13g2_fill_1
XFILLER_81_546 VPWR VGND sg13g2_fill_2
XFILLER_81_524 VPWR VGND sg13g2_fill_1
XFILLER_53_226 VPWR VGND sg13g2_fill_2
XFILLER_35_930 VPWR VGND sg13g2_fill_1
XFILLER_50_911 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2435 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1
+ VPWR i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[473\] clknet_leaf_114_clk sg13g2_dfrbpq_1
Xhold820 i_snitch.i_snitch_regfile.mem\[138\] VPWR VGND net852 sg13g2_dlygate4sd3_1
Xhold842 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold864 i_snitch.i_snitch_regfile.mem\[235\] VPWR VGND net896 sg13g2_dlygate4sd3_1
Xhold831 i_snitch.i_snitch_regfile.mem\[211\] VPWR VGND net863 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold853 i_snitch.i_snitch_regfile.mem\[199\] VPWR VGND net885 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2325 net1150 net2899 net2893 VPWR VGND sg13g2_a22oi_1
XFILLER_104_935 VPWR VGND sg13g2_decap_8
XFILLER_89_635 VPWR VGND sg13g2_fill_1
Xhold875 rsp_data_q\[20\] VPWR VGND net907 sg13g2_dlygate4sd3_1
Xhold897 i_snitch.i_snitch_regfile.mem\[83\] VPWR VGND net929 sg13g2_dlygate4sd3_1
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
Xhold886 i_snitch.i_snitch_regfile.mem\[230\] VPWR VGND net918 sg13g2_dlygate4sd3_1
XFILLER_77_808 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2471 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ net93 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_85_885 VPWR VGND sg13g2_decap_8
XFILLER_72_502 VPWR VGND sg13g2_decap_4
XFILLER_17_407 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N
+ VGND net3145 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N
+ sg13g2_o21ai_1
XFILLER_44_237 VPWR VGND sg13g2_fill_1
XFILLER_38_790 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1
+ net1400 VPWR VGND sg13g2_inv_2
XFILLER_26_963 VPWR VGND sg13g2_decap_8
XFILLER_73_1015 VPWR VGND sg13g2_decap_8
Xi_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_nand2_2
XFILLER_53_771 VPWR VGND sg13g2_fill_2
XFILLER_26_996 VPWR VGND sg13g2_fill_1
XFILLER_41_911 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2703 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2615 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2298 net1051 net2494 net1252 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[15\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net967 data_pdata\[15\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
Xstrb_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2729 strb_reg_q\[5\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D strb_reg_q\[4\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_12_112 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ net2561 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
XFILLER_8_149 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2887
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_294 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2576 net61 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B
+ net2564 sg13g2_a21oi_1
XFILLER_80_1008 VPWR VGND sg13g2_decap_8
XFILLER_79_145 VPWR VGND sg13g2_fill_2
XFILLER_79_134 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2716 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_67_318 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y net2840 i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_0_583 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[7\]
+ VGND net2293 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_48_565 VPWR VGND sg13g2_decap_8
XFILLER_36_705 VPWR VGND sg13g2_fill_1
XFILLER_91_877 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_440 VPWR VGND sg13g2_fill_2
XFILLER_73_70 VPWR VGND sg13g2_fill_2
XFILLER_16_473 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y net2637
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[493\] clknet_leaf_88_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_a22oi_1_B2_Y
+ net2323 net683 net2433 net2254 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2467 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_2
XFILLER_89_1000 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0 net3005 i_snitch.i_snitch_regfile.mem\[284\]
+ i_snitch.i_snitch_regfile.mem\[316\] i_snitch.i_snitch_regfile.mem\[348\] i_snitch.i_snitch_regfile.mem\[380\]
+ net2977 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2818 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND net2584 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[66\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[66\]
+ i_snitch.i_snitch_regfile.mem\[98\] net3117 i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_99_944 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_101_938 VPWR VGND sg13g2_decap_8
XFILLER_67_841 VPWR VGND sg13g2_fill_1
XFILLER_39_521 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR net916 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2463
+ net2254 net2659 net2860 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[65\] VGND sg13g2_inv_1
XFILLER_27_716 VPWR VGND sg13g2_decap_8
XFILLER_27_727 VPWR VGND sg13g2_fill_2
XFILLER_39_587 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A
+ VGND i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ sg13g2_o21ai_1
XFILLER_66_384 VPWR VGND sg13g2_decap_8
XFILLER_54_524 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VGND i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1
+ sg13g2_o21ai_1
XFILLER_82_888 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[316\] VGND sg13g2_inv_1
XFILLER_26_259 VPWR VGND sg13g2_decap_8
XFILLER_42_708 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[312\] clknet_leaf_67_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2958
+ i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2965
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_33_1021 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[337\] net2951 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0 net3137 i_snitch.i_snitch_regfile.mem\[408\]
+ i_snitch.i_snitch_regfile.mem\[440\] i_snitch.i_snitch_regfile.mem\[472\] i_snitch.i_snitch_regfile.mem\[504\]
+ net3111 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2538 sg13g2_a21oi_1
Xfanout2818 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y
+ net2818 VPWR VGND sg13g2_buf_8
Xhold650 data_pdata\[7\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net682 sg13g2_dlygate4sd3_1
Xfanout2807 net2808 net2807 VPWR VGND sg13g2_buf_8
Xhold672 i_snitch.i_snitch_regfile.mem\[269\] VPWR VGND net704 sg13g2_dlygate4sd3_1
Xhold661 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y VPWR VGND net693 sg13g2_dlygate4sd3_1
XFILLER_103_231 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_C
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X
+ VPWR VGND sg13g2_or4_1
Xhold683 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\] VPWR
+ VGND net715 sg13g2_dlygate4sd3_1
XFILLER_2_859 VPWR VGND sg13g2_decap_8
Xhold694 data_pdata\[13\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net726 sg13g2_dlygate4sd3_1
Xfanout2829 net2830 net2829 VPWR VGND sg13g2_buf_8
XFILLER_89_498 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y
+ sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[29\] net777 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_94_14 VPWR VGND sg13g2_decap_8
XFILLER_92_619 VPWR VGND sg13g2_fill_2
Xhold1350 rsp_data_q\[1\] VPWR VGND net1382 sg13g2_dlygate4sd3_1
Xhold1361 i_req_arb.data_i\[39\] VPWR VGND net1393 sg13g2_dlygate4sd3_1
XFILLER_57_340 VPWR VGND sg13g2_fill_2
XFILLER_85_693 VPWR VGND sg13g2_decap_4
Xhold1372 i_snitch.i_snitch_lsu.metadata_q\[2\] VPWR VGND net1404 sg13g2_dlygate4sd3_1
XFILLER_17_215 VPWR VGND sg13g2_decap_4
XFILLER_18_749 VPWR VGND sg13g2_decap_8
XFILLER_73_888 VPWR VGND sg13g2_fill_2
Xdata_pdata\[31\]_sg13g2_mux2_1_A1 rsp_data_q\[31\] net858 net3050 data_pdata\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_60_505 VPWR VGND sg13g2_fill_1
XFILLER_45_579 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[8\]_sg13g2_a22oi_1_A1 shift_reg_q\[8\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1_X
+ net3057 net3047 shift_reg_q\[8\] VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_25_292 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2321
+ sg13g2_o21ai_1
XFILLER_9_447 VPWR VGND sg13g2_fill_1
XFILLER_13_498 VPWR VGND sg13g2_decap_4
XFILLER_5_642 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[437\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2463 net2268 net2384 net1296 VPWR VGND sg13g2_a22oi_1
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_96_936 VPWR VGND sg13g2_decap_8
XFILLER_95_402 VPWR VGND sg13g2_decap_8
XFILLER_1_881 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q net3308 VGND VPWR i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[332\] clknet_leaf_71_clk sg13g2_dfrbpq_1
XFILLER_83_608 VPWR VGND sg13g2_decap_8
XFILLER_49_863 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[121\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[121\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2448 net2267 net2409 net1172 VPWR VGND sg13g2_a22oi_1
XFILLER_48_373 VPWR VGND sg13g2_fill_1
XFILLER_63_332 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[41\]
+ net2982 sg13g2_o21ai_1
XFILLER_51_505 VPWR VGND sg13g2_fill_1
XFILLER_36_546 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_or4_1_X
+ net3104 net3125 net3089 net3093 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B
+ VPWR VGND sg13g2_or4_1
XFILLER_16_281 VPWR VGND sg13g2_decap_4
XFILLER_104_1019 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[20\]_sg13g2_a22oi_1_A1 shift_reg_q\[20\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1_X
+ net3057 net3047 net496 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2379
+ sg13g2_o21ai_1
XFILLER_9_992 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_o21ai_1_A2
+ net3054 VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ VGND net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net104 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
XFILLER_98_240 VPWR VGND sg13g2_decap_4
XFILLER_101_702 VPWR VGND sg13g2_fill_2
XFILLER_98_273 VPWR VGND sg13g2_decap_8
XFILLER_101_746 VPWR VGND sg13g2_decap_8
XFILLER_100_212 VPWR VGND sg13g2_decap_8
XFILLER_87_958 VPWR VGND sg13g2_decap_8
XFILLER_104_35 VPWR VGND sg13g2_decap_8
XFILLER_95_980 VPWR VGND sg13g2_decap_8
XFILLER_100_289 VPWR VGND sg13g2_decap_8
XFILLER_55_822 VPWR VGND sg13g2_decap_4
XFILLER_39_395 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_93_clk clknet_5_20__leaf_clk clknet_leaf_93_clk VPWR VGND sg13g2_buf_8
XFILLER_15_708 VPWR VGND sg13g2_fill_2
XFILLER_70_847 VPWR VGND sg13g2_decap_4
XFILLER_70_836 VPWR VGND sg13g2_decap_4
XFILLER_42_549 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_a21o_1_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1 net2527 VPWR VGND sg13g2_xnor2_1
XFILLER_70_1018 VPWR VGND sg13g2_decap_8
XFILLER_22_251 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[457\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2376 net788 net2685 net2740 VPWR VGND sg13g2_a22oi_1
XFILLER_10_424 VPWR VGND sg13g2_fill_2
XFILLER_13_43 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q net3255 VGND VPWR i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[352\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_6_428 VPWR VGND sg13g2_fill_2
Xfanout3305 net3306 net3305 VPWR VGND sg13g2_buf_8
Xfanout3327 net3328 net3327 VPWR VGND sg13g2_buf_8
Xfanout3316 net3326 net3316 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net959 net2689 net2889 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2825
+ sg13g2_a221oi_1
Xfanout2604 net2605 net2604 VPWR VGND sg13g2_buf_2
Xfanout2615 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C_Y
+ net2615 VPWR VGND sg13g2_buf_8
XFILLER_78_903 VPWR VGND sg13g2_fill_2
Xfanout2626 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X
+ net2626 VPWR VGND sg13g2_buf_8
Xhold480 shift_reg_q\[23\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net512 sg13g2_dlygate4sd3_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_656 VPWR VGND sg13g2_decap_8
Xfanout2637 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y
+ net2637 VPWR VGND sg13g2_buf_8
Xfanout2648 data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y net2648 VPWR
+ VGND sg13g2_buf_2
Xfanout2659 net2660 net2659 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_o21ai_1_A1 net3012 VPWR i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[61\] net2985 sg13g2_o21ai_1
Xhold491 i_snitch.i_snitch_regfile.mem\[80\] VPWR VGND net523 sg13g2_dlygate4sd3_1
XFILLER_49_115 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2399
+ sg13g2_o21ai_1
XFILLER_92_449 VPWR VGND sg13g2_fill_1
XFILLER_92_438 VPWR VGND sg13g2_fill_1
XFILLER_79_1021 VPWR VGND sg13g2_decap_8
XFILLER_58_671 VPWR VGND sg13g2_fill_1
XFILLER_45_321 VPWR VGND sg13g2_fill_1
Xhold1191 rsp_data_q\[11\] VPWR VGND net1223 sg13g2_dlygate4sd3_1
Xhold1180 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] VPWR
+ VGND net1212 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_84_clk clknet_5_23__leaf_clk clknet_leaf_84_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2815 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A
+ VPWR VGND sg13g2_and2_1
XFILLER_60_346 VPWR VGND sg13g2_fill_1
XFILLER_33_538 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_13_251 VPWR VGND sg13g2_fill_1
XFILLER_9_222 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[51\] VGND sg13g2_inv_1
Xi_snitch.inst_addr_o\[12\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.pc_d\[12\]
+ i_snitch.inst_addr_o\[12\] clknet_leaf_57_clk sg13g2_dfrbpq_2
XFILLER_70_60 VPWR VGND sg13g2_fill_1
Xclkload25 clkload25/Y clknet_leaf_47_clk VPWR VGND sg13g2_inv_2
Xclkload14 clkload14/Y clknet_leaf_15_clk VPWR VGND sg13g2_inv_2
XFILLER_9_288 VPWR VGND sg13g2_fill_1
XFILLER_86_1014 VPWR VGND sg13g2_decap_8
Xclkload58 VPWR clkload58/Y clknet_leaf_64_clk VGND sg13g2_inv_1
Xclkload47 clknet_leaf_83_clk clkload47/Y VPWR VGND sg13g2_inv_4
Xclkload36 clkload36/Y clknet_leaf_105_clk VPWR VGND sg13g2_inv_2
XFILLER_6_984 VPWR VGND sg13g2_decap_8
XFILLER_5_472 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2552 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ sg13g2_a21oi_1
XFILLER_96_788 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
XFILLER_68_479 VPWR VGND sg13g2_fill_2
XFILLER_37_800 VPWR VGND sg13g2_decap_4
XFILLER_77_991 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net932 net2461 net2250 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q
+ net3241 VGND VPWR net955 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2832
+ VPWR i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[480\]
+ net2802 i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_75_clk clknet_5_19__leaf_clk clknet_leaf_75_clk VPWR VGND sg13g2_buf_8
XFILLER_93_1007 VPWR VGND sg13g2_decap_8
XFILLER_92_983 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2_sg13g2_inv_1_Y VPWR
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2 i_snitch.inst_addr_o\[13\]
+ VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_52_836 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q net3316 VGND VPWR i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[372\] clknet_leaf_66_clk sg13g2_dfrbpq_1
XFILLER_52_869 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1 VPWR VGND net3100 net2821
+ i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[58\]
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y net2824 sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q
+ net3191 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
Xclkload8 clknet_leaf_11_clk clkload8/X VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2
+ VGND net2747 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ sg13g2_o21ai_1
XFILLER_105_315 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y
+ net2566 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_o21ai_1_A1 net2970 VPWR i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[368\] net2805 sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A
+ i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a21oi_1_A1_B1 net2930 net2938 VPWR VGND
+ sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ VPWR VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_nand2b_2
XFILLER_8_1025 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[507\] clknet_leaf_117_clk sg13g2_dfrbpq_1
XFILLER_87_788 VPWR VGND sg13g2_decap_8
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0
+ net1122 i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y net2512
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_27_310 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y
+ net2611 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_66_clk clknet_5_27__leaf_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[49\] clknet_leaf_82_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_24_97 VPWR VGND sg13g2_fill_1
XFILLER_6_214 VPWR VGND sg13g2_fill_2
XFILLER_6_258 VPWR VGND sg13g2_fill_2
XFILLER_40_30 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C_sg13g2_inv_1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C
+ VGND sg13g2_inv_1
Xfanout3113 net3114 net3113 VPWR VGND sg13g2_buf_8
Xfanout3102 net3105 net3102 VPWR VGND sg13g2_buf_8
Xfanout3146 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_X
+ net3146 VPWR VGND sg13g2_buf_8
Xfanout3124 net3125 net3124 VPWR VGND sg13g2_buf_8
Xfanout3135 net3139 net3135 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[497\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net956 net2664 net2859 VPWR VGND sg13g2_a22oi_1
XFILLER_6_0 VPWR VGND sg13g2_decap_8
Xfanout2401 net2406 net2401 VPWR VGND sg13g2_buf_8
XFILLER_105_882 VPWR VGND sg13g2_decap_8
Xfanout3179 net3180 net3179 VPWR VGND sg13g2_buf_8
Xfanout2412 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y
+ net2412 VPWR VGND sg13g2_buf_8
XFILLER_3_976 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_fill_2
Xfanout3168 net3173 net3168 VPWR VGND sg13g2_buf_8
Xfanout2434 net2435 net2434 VPWR VGND sg13g2_buf_8
Xfanout2423 net2428 net2423 VPWR VGND sg13g2_buf_8
Xfanout3157 net3158 net3157 VPWR VGND sg13g2_buf_2
XFILLER_104_392 VPWR VGND sg13g2_decap_8
Xfanout2467 net2468 net2467 VPWR VGND sg13g2_buf_8
Xfanout2456 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y net2456 VPWR
+ VGND sg13g2_buf_8
Xfanout2445 net2447 net2445 VPWR VGND sg13g2_buf_8
Xfanout2478 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2478 VPWR VGND sg13g2_buf_8
XFILLER_78_766 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2340
+ sg13g2_o21ai_1
Xfanout2489 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y
+ net2489 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[392\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_93_736 VPWR VGND sg13g2_fill_2
XFILLER_65_416 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
XFILLER_59_980 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[181\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[181\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2443 net2268 net2342 net1175 VPWR VGND sg13g2_a22oi_1
XFILLER_1_35 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3094 i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
Xclkbuf_leaf_57_clk clknet_5_30__leaf_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
XFILLER_46_652 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2463 net2865 i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_18_376 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_33_324 VPWR VGND sg13g2_fill_2
XFILLER_61_688 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ net2611 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1
+ net2753 net3133 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_53_1024 VPWR VGND sg13g2_decap_4
XFILLER_14_593 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2782
+ i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2538 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2572 sg13g2_a21oi_2
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y net711 VPWR i_snitch.sb_d\[14\] VGND net2293
+ i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_and4_1_X
+ net3033 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C
+ VPWR VGND sg13g2_and4_1
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2431 net2247 net2317 net1171 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[69\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[69\] clknet_leaf_112_clk sg13g2_dfrbpq_1
XFILLER_102_329 VPWR VGND sg13g2_decap_8
XFILLER_68_221 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[211\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2542 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1
+ net47 sg13g2_a21oi_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.inst_addr_o\[21\] net2526 VPWR VGND sg13g2_nand2_1
XFILLER_60_1028 VPWR VGND sg13g2_fill_1
Xfanout2990 net2995 net2990 VPWR VGND sg13g2_buf_8
XFILLER_68_298 VPWR VGND sg13g2_fill_2
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X net2480 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X
+ net2498 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_48_clk clknet_5_13__leaf_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C
+ net2710 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C_Y
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.i_snitch_regfile.mem\[317\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[317\]
+ net3012 i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_a21oi_1_A1_Y net2985 sg13g2_a21oi_1
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_37_685 VPWR VGND sg13g2_fill_1
XFILLER_101_14 VPWR VGND sg13g2_decap_8
XFILLER_80_931 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2846
+ sg13g2_a221oi_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2
+ net2506 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_40_806 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net2555 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
XFILLER_106_624 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_105_112 VPWR VGND sg13g2_decap_8
XFILLER_79_519 VPWR VGND sg13g2_decap_4
XFILLER_105_189 VPWR VGND sg13g2_decap_8
XFILLER_102_863 VPWR VGND sg13g2_decap_8
XFILLER_86_59 VPWR VGND sg13g2_fill_2
XFILLER_48_906 VPWR VGND sg13g2_decap_4
XFILLER_0_968 VPWR VGND sg13g2_decap_8
XFILLER_47_416 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_39_clk clknet_5_10__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_75_758 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B VPWR
+ VGND sg13g2_nor2_1
XFILLER_28_652 VPWR VGND sg13g2_fill_2
XFILLER_56_983 VPWR VGND sg13g2_decap_4
XFILLER_55_471 VPWR VGND sg13g2_decap_8
XFILLER_55_482 VPWR VGND sg13g2_fill_1
XFILLER_15_346 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]
+ net3176 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_71_997 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[270\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q net3215 VGND VPWR i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[89\] clknet_leaf_113_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ net2593 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[231\] clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_100_1022 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_B_N i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2
+ VPWR VGND sg13g2_nor2b_1
XFILLER_83_1028 VPWR VGND sg13g2_fill_1
Xfanout2242 net2243 net2242 VPWR VGND sg13g2_buf_8
Xfanout2253 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2253 VPWR VGND sg13g2_buf_8
Xdata_pdata\[10\]_sg13g2_nor2b_1_A data_pdata\[10\] net3157 data_pdata\[10\]_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
Xfanout2264 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ net2264 VPWR VGND sg13g2_buf_8
Xfanout2286 net2287 net2286 VPWR VGND sg13g2_buf_8
Xfanout2275 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2275 VPWR VGND sg13g2_buf_8
Xfanout2297 net2298 net2297 VPWR VGND sg13g2_buf_8
XFILLER_93_544 VPWR VGND sg13g2_fill_2
XFILLER_65_268 VPWR VGND sg13g2_fill_2
XFILLER_46_471 VPWR VGND sg13g2_fill_1
XFILLER_34_644 VPWR VGND sg13g2_decap_4
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X VGND
+ VPWR i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2 i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C
+ sg13g2_or2_1
XFILLER_21_338 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2632 VPWR i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xshift_reg_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2735 shift_reg_q\[20\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[16\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[16\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_89_839 VPWR VGND sg13g2_decap_8
XFILLER_88_316 VPWR VGND sg13g2_fill_2
XFILLER_0_209 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_nor3_1_A net1370 net2885 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_102_126 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_97_894 VPWR VGND sg13g2_decap_8
XFILLER_96_382 VPWR VGND sg13g2_fill_2
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_449 VPWR VGND sg13g2_decap_4
XFILLER_53_920 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ VGND i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y
+ net33 sg13g2_o21ai_1
XFILLER_53_975 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[251\] clknet_leaf_119_clk sg13g2_dfrbpq_1
XFILLER_24_121 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[70\]
+ net2846 i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
XFILLER_21_850 VPWR VGND sg13g2_fill_2
XFILLER_97_14 VPWR VGND sg13g2_decap_8
XFILLER_4_537 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_or2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2
+ net2924 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1
+ sg13g2_a21oi_1
XFILLER_88_861 VPWR VGND sg13g2_decap_8
XFILLER_0_765 VPWR VGND sg13g2_decap_8
XFILLER_94_319 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ net2545 net2703 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_87_360 VPWR VGND sg13g2_fill_1
XFILLER_75_500 VPWR VGND sg13g2_decap_8
XFILLER_48_758 VPWR VGND sg13g2_fill_2
XFILLER_90_503 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 net2755
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_547 VPWR VGND sg13g2_fill_2
XFILLER_43_474 VPWR VGND sg13g2_fill_1
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q
+ net3231 VGND VPWR net654 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_30_179 VPWR VGND sg13g2_fill_1
XFILLER_7_67 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[376\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2397 net1191 net2666 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_98_647 VPWR VGND sg13g2_fill_1
XFILLER_79_850 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[90\]
+ net2840 i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2870
+ net2676 VPWR VGND sg13g2_nand2_1
XFILLER_100_619 VPWR VGND sg13g2_decap_8
XFILLER_87_80 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[271\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xhold1009 i_snitch.i_snitch_regfile.mem\[205\] VPWR VGND net1041 sg13g2_dlygate4sd3_1
XFILLER_93_330 VPWR VGND sg13g2_fill_1
XFILLER_16_2 VPWR VGND sg13g2_fill_1
XFILLER_38_246 VPWR VGND sg13g2_fill_1
XFILLER_94_875 VPWR VGND sg13g2_decap_8
XFILLER_93_352 VPWR VGND sg13g2_fill_2
XFILLER_66_588 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[377\]
+ net3119 i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_a21oi_1_A1_Y net2941 sg13g2_a21oi_1
XFILLER_62_794 VPWR VGND sg13g2_fill_1
XFILLER_62_772 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2788
+ net2659 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y net3129 sg13g2_o21ai_1
XFILLER_34_463 VPWR VGND sg13g2_fill_2
XFILLER_34_496 VPWR VGND sg13g2_fill_1
XFILLER_50_989 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q net3316 VGND VPWR i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[406\] clknet_leaf_65_clk sg13g2_dfrbpq_2
XFILLER_30_680 VPWR VGND sg13g2_fill_1
Xhold821 i_snitch.i_snitch_regfile.mem\[150\] VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold810 i_snitch.i_snitch_regfile.mem\[511\] VPWR VGND net842 sg13g2_dlygate4sd3_1
XFILLER_104_914 VPWR VGND sg13g2_decap_8
XFILLER_66_1023 VPWR VGND sg13g2_decap_4
Xhold832 i_snitch.i_snitch_regfile.mem\[340\] VPWR VGND net864 sg13g2_dlygate4sd3_1
Xhold854 i_snitch.i_snitch_regfile.mem\[416\] VPWR VGND net886 sg13g2_dlygate4sd3_1
Xhold843 i_snitch.i_snitch_regfile.mem\[489\] VPWR VGND net875 sg13g2_dlygate4sd3_1
XFILLER_103_413 VPWR VGND sg13g2_fill_2
Xhold876 rsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net908 sg13g2_dlygate4sd3_1
Xhold865 i_snitch.i_snitch_regfile.mem\[171\] VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold898 i_snitch.i_snitch_regfile.mem\[362\] VPWR VGND net930 sg13g2_dlygate4sd3_1
Xhold887 i_snitch.i_snitch_regfile.mem\[74\] VPWR VGND net919 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_A1
+ VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ sg13g2_or2_1
XFILLER_97_680 VPWR VGND sg13g2_decap_8
XFILLER_88_179 VPWR VGND sg13g2_fill_2
XFILLER_69_360 VPWR VGND sg13g2_fill_1
XFILLER_85_864 VPWR VGND sg13g2_decap_8
XFILLER_84_363 VPWR VGND sg13g2_fill_1
XFILLER_45_728 VPWR VGND sg13g2_decap_4
XFILLER_45_706 VPWR VGND sg13g2_decap_8
XFILLER_29_246 VPWR VGND sg13g2_fill_1
Xcnt_q\[0\]_sg13g2_dfrbpq_1_Q net3184 VGND VPWR cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D cnt_q\[0\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_2
XFILLER_53_750 VPWR VGND sg13g2_fill_1
XFILLER_80_580 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y net2518
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 VPWR VGND sg13g2_inv_4
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net1121 net2691 net3041 VPWR VGND sg13g2_a22oi_1
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_32_75 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[291\] clknet_leaf_104_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2480 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2498 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_0 VPWR VGND sg13g2_decap_8
XFILLER_106_273 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xrsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ net908 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2872
+ net2661 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y sg13g2_or2_1
XFILLER_103_991 VPWR VGND sg13g2_decap_8
XFILLER_63_503 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2431
+ net2275 VPWR VGND sg13g2_nand2_1
XFILLER_91_856 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_430 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[426\] clknet_leaf_101_clk sg13g2_dfrbpq_1
XFILLER_35_249 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[215\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net791 net2648 net2791 VPWR VGND sg13g2_a22oi_1
XFILLER_32_945 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[110\] clknet_leaf_83_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0 net3006 i_snitch.i_snitch_regfile.mem\[131\]
+ i_snitch.i_snitch_regfile.mem\[163\] i_snitch.i_snitch_regfile.mem\[195\] i_snitch.i_snitch_regfile.mem\[227\]
+ net2979 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_99_923 VPWR VGND sg13g2_decap_8
XFILLER_98_422 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1049 net708 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_101_917 VPWR VGND sg13g2_decap_8
XFILLER_98_499 VPWR VGND sg13g2_fill_1
XFILLER_86_617 VPWR VGND sg13g2_decap_8
XFILLER_79_680 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C
+ net2756 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_58_319 VPWR VGND sg13g2_decap_8
XFILLER_100_427 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2774
+ net2668 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2640 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_66_363 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[106\]
+ net2804 sg13g2_o21ai_1
XFILLER_96_1027 VPWR VGND sg13g2_fill_2
XFILLER_82_867 VPWR VGND sg13g2_decap_8
XFILLER_81_344 VPWR VGND sg13g2_decap_8
XFILLER_26_238 VPWR VGND sg13g2_decap_8
XFILLER_22_433 VPWR VGND sg13g2_fill_2
XFILLER_23_945 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A_Y net2845 i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2399
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1343 net2491 net1377 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[24\] net712 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_50_797 VPWR VGND sg13g2_fill_1
XFILLER_10_639 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A_sg13g2_nand3_1_Y
+ net3073 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B
+ net3034 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A
+ VPWR VGND sg13g2_nand3_1
XFILLER_5_109 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[42\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2474 VPWR VGND sg13g2_nand2_1
Xhold651 i_snitch.i_snitch_regfile.mem\[282\] VPWR VGND net683 sg13g2_dlygate4sd3_1
XFILLER_2_838 VPWR VGND sg13g2_decap_8
Xhold640 i_snitch.i_snitch_regfile.mem\[338\] VPWR VGND net672 sg13g2_dlygate4sd3_1
Xhold662 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y VPWR VGND net694 sg13g2_dlygate4sd3_1
Xfanout2819 net2820 net2819 VPWR VGND sg13g2_buf_8
Xfanout2808 net2809 net2808 VPWR VGND sg13g2_buf_8
XFILLER_103_210 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2
+ VPWR VGND sg13g2_nor3_1
Xhold673 i_snitch.i_snitch_regfile.mem\[172\] VPWR VGND net705 sg13g2_dlygate4sd3_1
Xhold684 i_snitch.i_snitch_regfile.mem\[471\] VPWR VGND net716 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2642 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xhold695 i_snitch.i_snitch_regfile.mem\[177\] VPWR VGND net727 sg13g2_dlygate4sd3_1
XFILLER_104_788 VPWR VGND sg13g2_decap_8
XFILLER_77_628 VPWR VGND sg13g2_fill_2
XFILLER_49_319 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[446\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_103_287 VPWR VGND sg13g2_decap_8
XFILLER_76_138 VPWR VGND sg13g2_fill_1
Xhold1340 i_snitch.inst_addr_o\[23\] VPWR VGND net1372 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[235\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[235\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net896 net2679 net2875 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2861
+ net2669 VPWR VGND sg13g2_nand2_1
Xhold1351 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] VPWR
+ VGND net1383 sg13g2_dlygate4sd3_1
XFILLER_40_1026 VPWR VGND sg13g2_fill_2
XFILLER_100_994 VPWR VGND sg13g2_decap_8
Xhold1362 i_snitch.inst_addr_o\[20\] VPWR VGND net1394 sg13g2_dlygate4sd3_1
Xhold1373 i_req_arb.data_i\[43\] VPWR VGND net1405 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[275\] VGND sg13g2_inv_1
XFILLER_18_728 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ net2584 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[130\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_72_388 VPWR VGND sg13g2_fill_2
XFILLER_60_517 VPWR VGND sg13g2_fill_1
XFILLER_14_912 VPWR VGND sg13g2_decap_8
XFILLER_26_783 VPWR VGND sg13g2_fill_2
XFILLER_14_967 VPWR VGND sg13g2_fill_1
XFILLER_41_731 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_nand2_1_A_Y net3029 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A_Y VPWR VGND sg13g2_a22oi_1
XFILLER_43_74 VPWR VGND sg13g2_decap_8
XFILLER_9_415 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y net3012 sg13g2_o21ai_1
XFILLER_40_285 VPWR VGND sg13g2_fill_1
XFILLER_41_797 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2489 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ sg13g2_o21ai_1
XFILLER_5_621 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_96_915 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2549 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_68_628 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[341\] net2948 VPWR VGND sg13g2_nand2_1
XFILLER_1_860 VPWR VGND sg13g2_decap_8
XFILLER_95_436 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[27\]_sg13g2_dfrbpq_1_Q net3238 VGND VPWR rsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[27\] clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_49_875 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0 net3126 i_snitch.i_snitch_regfile.mem\[412\]
+ i_snitch.i_snitch_regfile.mem\[444\] i_snitch.i_snitch_regfile.mem\[476\] i_snitch.i_snitch_regfile.mem\[508\]
+ net3106 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_90_130 VPWR VGND sg13g2_fill_2
XFILLER_36_569 VPWR VGND sg13g2_decap_8
XFILLER_63_366 VPWR VGND sg13g2_fill_2
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2_1_B
+ i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_16_260 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_937 VPWR VGND sg13g2_fill_2
XFILLER_69_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[466\] clknet_leaf_90_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[255\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2330 net761 net2646 net2874 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2610 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_99_797 VPWR VGND sg13g2_decap_8
XFILLER_87_937 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[150\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_86_436 VPWR VGND sg13g2_fill_2
XFILLER_104_14 VPWR VGND sg13g2_decap_8
XFILLER_100_268 VPWR VGND sg13g2_decap_8
XFILLER_39_352 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2920
+ sg13g2_a221oi_1
Xi_req_arb.data_i\[41\]_sg13g2_inv_1_A i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_A1 net1361
+ VPWR VGND sg13g2_inv_2
XFILLER_66_193 VPWR VGND sg13g2_decap_8
XFILLER_70_815 VPWR VGND sg13g2_fill_1
XFILLER_23_742 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2720 i_snitch.inst_addr_o\[27\] sg13g2_a21oi_2
XFILLER_7_908 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2578 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xshift_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2736 shift_reg_q\[8\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[4\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2436 net2872 i_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q_D net2905
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2607 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2364
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ net3026 net2974 VPWR VGND sg13g2_nand2_2
Xfanout3328 net3329 net3328 VPWR VGND sg13g2_buf_8
Xfanout3317 net3326 net3317 VPWR VGND sg13g2_buf_8
Xfanout3306 net3313 net3306 VPWR VGND sg13g2_buf_8
Xfanout2605 net2606 net2605 VPWR VGND sg13g2_buf_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A
+ net3145 VPWR VGND net3142 sg13g2_nand2b_2
Xfanout2627 net2628 net2627 VPWR VGND sg13g2_buf_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_2_635 VPWR VGND sg13g2_decap_8
Xhold470 strb_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold481 i_snitch.i_snitch_regfile.mem\[458\] VPWR VGND net513 sg13g2_dlygate4sd3_1
Xfanout2616 net2618 net2616 VPWR VGND sg13g2_buf_8
XFILLER_104_563 VPWR VGND sg13g2_decap_8
Xfanout2649 net2650 net2649 VPWR VGND sg13g2_buf_8
Xfanout2638 net2640 net2638 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0 net3128 i_snitch.i_snitch_regfile.mem\[138\]
+ i_snitch.i_snitch_regfile.mem\[170\] i_snitch.i_snitch_regfile.mem\[202\] i_snitch.i_snitch_regfile.mem\[234\]
+ net3107 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold492 i_snitch.i_snitch_regfile.mem\[417\] VPWR VGND net524 sg13g2_dlygate4sd3_1
XFILLER_78_959 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.inst_addr_o\[23\] net2525 VPWR VGND sg13g2_xnor2_1
XFILLER_38_30 VPWR VGND sg13g2_fill_2
XFILLER_79_1000 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2b_1
XFILLER_57_171 VPWR VGND sg13g2_fill_1
Xhold1170 i_snitch.i_snitch_regfile.mem\[444\] VPWR VGND net1202 sg13g2_dlygate4sd3_1
XFILLER_18_525 VPWR VGND sg13g2_fill_2
XFILLER_100_791 VPWR VGND sg13g2_decap_8
Xhold1192 rsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1224
+ sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2854
+ net2674 VPWR VGND sg13g2_nand2_1
Xhold1181 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] VPWR
+ VGND net1213 sg13g2_dlygate4sd3_1
XFILLER_61_837 VPWR VGND sg13g2_decap_8
XFILLER_45_366 VPWR VGND sg13g2_fill_2
XFILLER_72_174 VPWR VGND sg13g2_fill_2
XFILLER_61_848 VPWR VGND sg13g2_fill_1
Xdata_pdata\[29\]_sg13g2_nand2b_1_B data_pdata\[29\]_sg13g2_nand2b_1_B_Y data_pdata\[29\]
+ net3155 VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[486\] clknet_leaf_77_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q_D VGND net2315 net310
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2323 net1143 net2433 net2270 VPWR VGND sg13g2_a22oi_1
XFILLER_9_201 VPWR VGND sg13g2_decap_8
XFILLER_41_572 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_C
+ VPWR VGND sg13g2_nor4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2500 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xclkload26 VPWR clkload26/Y clknet_leaf_48_clk VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2818 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xclkload15 clknet_leaf_19_clk clkload15/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q net3278 VGND VPWR i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[170\] clknet_leaf_94_clk sg13g2_dfrbpq_1
Xclkload48 VPWR clkload48/Y clknet_leaf_50_clk VGND sg13g2_inv_1
Xclkload59 clknet_leaf_80_clk clkload59/X VPWR VGND sg13g2_buf_8
XFILLER_6_963 VPWR VGND sg13g2_decap_8
Xclkload37 clknet_leaf_75_clk clkload37/X VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nand2b_1_B i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C VPWR VGND net2867 sg13g2_nand2b_2
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_5_495 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[276\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[276\]
+ net3030 i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_a21oi_1_A1_Y net2993 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0 net3013 i_snitch.i_snitch_regfile.mem\[257\]
+ i_snitch.i_snitch_regfile.mem\[289\] i_snitch.i_snitch_regfile.mem\[385\] i_snitch.i_snitch_regfile.mem\[417\]
+ net2963 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_96_734 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VGND net2557 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ sg13g2_o21ai_1
XFILLER_96_778 VPWR VGND sg13g2_fill_1
Xdata_pdata\[28\]_sg13g2_dfrbpq_1_Q net3236 VGND VPWR data_pdata\[28\]_sg13g2_dfrbpq_1_Q_D
+ data_pdata\[28\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_48_160 VPWR VGND sg13g2_decap_8
XFILLER_92_962 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X
+ net2752 net2849 sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[305\] clknet_leaf_79_clk sg13g2_dfrbpq_1
XFILLER_36_355 VPWR VGND sg13g2_fill_1
XFILLER_52_848 VPWR VGND sg13g2_fill_1
XFILLER_17_580 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[77\]
+ i_snitch.i_snitch_regfile.mem\[109\] net3131 i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_51_358 VPWR VGND sg13g2_fill_2
XFILLER_20_745 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[261\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2478 i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2472 net2795 i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
Xclkload9 VPWR clkload9/Y clknet_leaf_12_clk VGND sg13g2_inv_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B sg13g2_o21ai_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ net2602 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_and2_1
XFILLER_99_572 VPWR VGND sg13g2_fill_2
XFILLER_8_1004 VPWR VGND sg13g2_decap_8
XFILLER_59_425 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_nand2b_1_A_N_Y
+ net3026 i_snitch.i_snitch_regfile.mem\[92\] VPWR VGND sg13g2_nand2b_1
XFILLER_87_778 VPWR VGND sg13g2_decap_4
XFILLER_75_907 VPWR VGND sg13g2_decap_4
XFILLER_74_439 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[348\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[348\] net2950 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[295\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2430 net2285 net2316 net1218 VPWR VGND sg13g2_a22oi_1
XFILLER_83_984 VPWR VGND sg13g2_decap_8
XFILLER_27_366 VPWR VGND sg13g2_fill_1
XFILLER_42_303 VPWR VGND sg13g2_fill_1
XFILLER_82_494 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[190\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_42_347 VPWR VGND sg13g2_decap_8
XFILLER_42_358 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[296\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[296\]
+ net3019 i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_a21oi_1_A1_Y net2990 sg13g2_a21oi_1
XFILLER_50_380 VPWR VGND sg13g2_fill_1
XFILLER_10_211 VPWR VGND sg13g2_decap_8
XFILLER_11_778 VPWR VGND sg13g2_fill_2
XFILLER_10_299 VPWR VGND sg13g2_fill_1
Xfanout3103 net3105 net3103 VPWR VGND sg13g2_buf_8
XFILLER_40_75 VPWR VGND sg13g2_fill_1
Xfanout3147 net3148 net3147 VPWR VGND sg13g2_buf_8
Xfanout3114 net3114 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_buf_16
Xfanout3136 net3139 net3136 VPWR VGND sg13g2_buf_8
Xfanout3125 net80 net3125 VPWR VGND sg13g2_buf_8
XFILLER_3_955 VPWR VGND sg13g2_decap_8
Xfanout2402 net2406 net2402 VPWR VGND sg13g2_buf_8
XFILLER_105_861 VPWR VGND sg13g2_decap_8
Xfanout3169 net3171 net3169 VPWR VGND sg13g2_buf_8
Xfanout2424 net2428 net2424 VPWR VGND sg13g2_buf_8
Xfanout2435 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2435 VPWR
+ VGND sg13g2_buf_8
Xfanout2413 i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ net2413 VPWR VGND sg13g2_buf_8
Xfanout3158 i_snitch.i_snitch_lsu.metadata_q\[2\] net3158 VPWR VGND sg13g2_buf_8
XFILLER_104_371 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor4_1_Y
+ net3077 net83 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2340
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[325\] clknet_leaf_110_clk sg13g2_dfrbpq_1
Xfanout2446 net2447 net2446 VPWR VGND sg13g2_buf_8
Xfanout2457 net2459 net2457 VPWR VGND sg13g2_buf_8
Xfanout2468 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2468 VPWR
+ VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_1_14 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2450 net2273 net2411 net1273 VPWR VGND sg13g2_a22oi_1
Xfanout2479 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y
+ net2479 VPWR VGND sg13g2_buf_8
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2855
+ i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_18_300 VPWR VGND sg13g2_decap_4
XFILLER_19_834 VPWR VGND sg13g2_fill_2
XFILLER_74_940 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2572 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2538 sg13g2_a21oi_1
XFILLER_74_984 VPWR VGND sg13g2_fill_2
XFILLER_73_472 VPWR VGND sg13g2_decap_4
XFILLER_46_664 VPWR VGND sg13g2_fill_2
XFILLER_45_196 VPWR VGND sg13g2_fill_1
XFILLER_60_177 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[13\]_sg13g2_a22oi_1_A1 shift_reg_q\[13\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ net3053 net3043 net476 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[391\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_A
+ VPWR i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1_A1 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_6_782 VPWR VGND sg13g2_fill_1
XFILLER_103_809 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B
+ VGND net2540 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A VPWR
+ VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y net3006 sg13g2_o21ai_1
XFILLER_102_308 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_88_509 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y
+ net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_69_756 VPWR VGND sg13g2_decap_4
Xfanout2991 net2995 net2991 VPWR VGND sg13g2_buf_8
Xfanout2980 net2984 net2980 VPWR VGND sg13g2_buf_8
XFILLER_69_789 VPWR VGND sg13g2_fill_2
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_84_759 VPWR VGND sg13g2_decap_4
XFILLER_37_642 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ net2744 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor4_1
XFILLER_80_910 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1
+ net1385 VPWR VGND sg13g2_inv_2
XFILLER_65_973 VPWR VGND sg13g2_fill_1
XFILLER_65_962 VPWR VGND sg13g2_decap_8
XFILLER_52_612 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net471 net2491 VPWR VGND sg13g2_nand2_1
XFILLER_80_987 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A
+ VPWR VGND sg13g2_nand2_2
XFILLER_52_678 VPWR VGND sg13g2_decap_4
XFILLER_20_531 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[345\] clknet_leaf_114_clk sg13g2_dfrbpq_1
XFILLER_20_553 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_106_614 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2350 net965 net2900 net2888 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_A1
+ net2307 i_snitch.pc_d\[24\] i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
XFILLER_106_669 VPWR VGND sg13g2_decap_8
XFILLER_105_168 VPWR VGND sg13g2_decap_8
XFILLER_87_520 VPWR VGND sg13g2_fill_1
XFILLER_0_947 VPWR VGND sg13g2_decap_8
XFILLER_102_842 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[0\]_sg13g2_nand2_1_Y i_snitch.pc_d\[0\] i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
XFILLER_59_244 VPWR VGND sg13g2_decap_8
XFILLER_59_233 VPWR VGND sg13g2_fill_2
Xi_snitch.gpr_waddr\[7\]_sg13g2_dfrbpq_1_Q net3251 VGND VPWR i_snitch.gpr_waddr\[7\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.gpr_waddr\[7\] clknet_leaf_19_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A_Y net2840 i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_101_385 VPWR VGND sg13g2_decap_4
XFILLER_90_729 VPWR VGND sg13g2_decap_8
XFILLER_90_718 VPWR VGND sg13g2_decap_8
XFILLER_76_1025 VPWR VGND sg13g2_decap_4
XFILLER_16_837 VPWR VGND sg13g2_fill_2
XFILLER_16_859 VPWR VGND sg13g2_fill_1
XFILLER_30_328 VPWR VGND sg13g2_fill_2
XFILLER_11_531 VPWR VGND sg13g2_decap_8
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_100_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_546 VPWR VGND sg13g2_fill_1
XFILLER_13_1020 VPWR VGND sg13g2_decap_8
XFILLER_7_568 VPWR VGND sg13g2_decap_8
XFILLER_98_829 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2
+ VPWR VGND net2924 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y
+ sg13g2_a221oi_1
XFILLER_3_752 VPWR VGND sg13g2_fill_2
Xfanout2243 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2243 VPWR VGND sg13g2_buf_8
Xfanout2276 net2277 net2276 VPWR VGND sg13g2_buf_8
Xfanout2265 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ net2265 VPWR VGND sg13g2_buf_8
Xfanout2254 net2255 net2254 VPWR VGND sg13g2_buf_8
XFILLER_25_7 VPWR VGND sg13g2_decap_4
Xdata_pdata\[3\]_sg13g2_mux2_1_A1 rsp_data_q\[3\] net688 net3048 data_pdata\[3\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_93_523 VPWR VGND sg13g2_fill_2
Xfanout2298 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_Y net2298 VPWR VGND
+ sg13g2_buf_8
XFILLER_65_214 VPWR VGND sg13g2_decap_8
Xfanout2287 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y
+ net2287 VPWR VGND sg13g2_buf_8
XFILLER_65_247 VPWR VGND sg13g2_fill_1
XFILLER_93_567 VPWR VGND sg13g2_decap_4
XFILLER_81_718 VPWR VGND sg13g2_fill_2
XFILLER_46_461 VPWR VGND sg13g2_fill_2
XFILLER_18_141 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1157 net3065 rsp_data_q\[26\] VPWR VGND sg13g2_a22oi_1
XFILLER_73_280 VPWR VGND sg13g2_fill_1
XFILLER_19_697 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q net3286 VGND VPWR i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[365\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_62_976 VPWR VGND sg13g2_decap_4
XFILLER_22_807 VPWR VGND sg13g2_fill_1
XFILLER_61_475 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net1009 net2445 net2254 VPWR VGND sg13g2_a22oi_1
XFILLER_30_840 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ VGND net2711 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_o21ai_1_A1 net3110 VPWR i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[74\] net3132 sg13g2_o21ai_1
XFILLER_89_818 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0
+ VGND net2606 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_103_639 VPWR VGND sg13g2_fill_1
XFILLER_102_105 VPWR VGND sg13g2_decap_8
XFILLER_99_1014 VPWR VGND sg13g2_decap_8
XFILLER_97_873 VPWR VGND sg13g2_decap_8
XFILLER_84_501 VPWR VGND sg13g2_fill_2
XFILLER_84_589 VPWR VGND sg13g2_fill_2
Xi_snitch.inst_addr_o\[25\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[25\]
+ i_snitch.inst_addr_o\[25\] clknet_leaf_52_clk sg13g2_dfrbpq_2
XFILLER_56_269 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2933 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
XFILLER_53_943 VPWR VGND sg13g2_decap_4
XFILLER_24_111 VPWR VGND sg13g2_fill_2
XFILLER_25_634 VPWR VGND sg13g2_decap_4
XFILLER_80_762 VPWR VGND sg13g2_decap_8
XFILLER_25_645 VPWR VGND sg13g2_fill_1
XFILLER_80_795 VPWR VGND sg13g2_fill_2
XFILLER_53_987 VPWR VGND sg13g2_fill_1
XFILLER_106_488 VPWR VGND sg13g2_decap_8
XFILLER_0_744 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q net3274 VGND VPWR i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[385\] clknet_leaf_103_clk sg13g2_dfrbpq_1
XFILLER_48_726 VPWR VGND sg13g2_fill_1
XFILLER_101_182 VPWR VGND sg13g2_decap_8
XFILLER_75_523 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[174\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2344 net974 net2688 net2774 VPWR VGND sg13g2_a22oi_1
XFILLER_29_940 VPWR VGND sg13g2_fill_2
XFILLER_44_943 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_71_751 VPWR VGND sg13g2_fill_1
XFILLER_102_91 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
XFILLER_31_615 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_15_188 VPWR VGND sg13g2_decap_8
XFILLER_11_350 VPWR VGND sg13g2_decap_8
XFILLER_12_873 VPWR VGND sg13g2_decap_4
XFILLER_7_46 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2432 net2269 net2316 net1221 VPWR VGND sg13g2_a22oi_1
XFILLER_98_615 VPWR VGND sg13g2_decap_8
XFILLER_98_604 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[204\] clknet_leaf_68_clk sg13g2_dfrbpq_1
XFILLER_94_854 VPWR VGND sg13g2_decap_8
XFILLER_38_236 VPWR VGND sg13g2_fill_1
XFILLER_54_729 VPWR VGND sg13g2_fill_2
XFILLER_81_548 VPWR VGND sg13g2_fill_1
XFILLER_81_537 VPWR VGND sg13g2_fill_1
XFILLER_62_740 VPWR VGND sg13g2_decap_4
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_19_494 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[266\] VGND sg13g2_inv_1
XFILLER_50_913 VPWR VGND sg13g2_fill_1
XFILLER_99_0 VPWR VGND sg13g2_decap_8
XFILLER_21_169 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_or2_1_A VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_or2_1_A_X
+ i_snitch.i_snitch_lsu.metadata_q\[1\] i_snitch.i_snitch_lsu.metadata_q\[0\] sg13g2_or2_1
Xhold800 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net832 sg13g2_dlygate4sd3_1
Xhold811 i_snitch.i_snitch_regfile.mem\[111\] VPWR VGND net843 sg13g2_dlygate4sd3_1
Xhold822 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\] VPWR
+ VGND net854 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[500\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2370 net969 net2671 net2857 VPWR VGND sg13g2_a22oi_1
Xhold833 i_snitch.i_snitch_regfile.mem\[256\] VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold855 i_snitch.i_snitch_regfile.mem\[155\] VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold844 i_snitch.i_snitch_regfile.mem\[94\] VPWR VGND net876 sg13g2_dlygate4sd3_1
Xhold888 i_snitch.i_snitch_regfile.mem\[56\] VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold866 i_snitch.i_snitch_regfile.mem\[407\] VPWR VGND net898 sg13g2_dlygate4sd3_1
Xhold877 i_snitch.i_snitch_regfile.mem\[348\] VPWR VGND net909 sg13g2_dlygate4sd3_1
XFILLER_88_147 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C
+ net2490 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nand3_1
Xhold899 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\] VPWR
+ VGND net931 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ net2697 net2541 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
XFILLER_85_843 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1168 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y net2282
+ VPWR VGND sg13g2_a22oi_1
XFILLER_53_773 VPWR VGND sg13g2_fill_1
XFILLER_52_261 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2402 net733 net2686 net2795 VPWR VGND sg13g2_a22oi_1
XFILLER_26_987 VPWR VGND sg13g2_fill_1
XFILLER_41_913 VPWR VGND sg13g2_fill_1
XFILLER_53_795 VPWR VGND sg13g2_fill_2
XFILLER_12_114 VPWR VGND sg13g2_fill_1
XFILLER_12_147 VPWR VGND sg13g2_decap_4
XFILLER_40_456 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[224\] clknet_leaf_49_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ net2544 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_q\[1\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[1\] i_snitch.sb_q\[1\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
Xstrb_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR strb_reg_q\[6\]_sg13g2_nand2_1_A_Y
+ strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A strb_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ strb_reg_q\[5\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[68\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2476 i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nor3_1_A_Y net2452 net2784 i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_dfrbpq_1_Q_D
+ net2908 sg13g2_a221oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C
+ net96 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_4_357 VPWR VGND sg13g2_decap_4
XFILLER_4_335 VPWR VGND sg13g2_decap_8
XFILLER_106_252 VPWR VGND sg13g2_decap_8
XFILLER_103_970 VPWR VGND sg13g2_decap_8
XFILLER_79_169 VPWR VGND sg13g2_fill_2
XFILLER_0_541 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2419 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_57_84 VPWR VGND sg13g2_decap_8
XFILLER_57_73 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_75_386 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1
+ i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_63_559 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X VPWR VGND
+ sg13g2_or3_1
XFILLER_17_965 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_92_7 VPWR VGND sg13g2_decap_8
XFILLER_32_935 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_692 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] net612 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_7_184 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_99_902 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1040 net2456 net2245 VPWR VGND sg13g2_a22oi_1
XFILLER_99_979 VPWR VGND sg13g2_decap_8
XFILLER_98_91 VPWR VGND sg13g2_decap_8
Xdata_pdata\[23\]_sg13g2_nor2b_1_B_N net3160 data_pdata\[23\] data_pdata\[23\]_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2405 net1073 net2473 net2251 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2636 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_B1
+ net669 net2301 VPWR VGND sg13g2_nand2_1
XFILLER_14_0 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2861
+ i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_96_1006 VPWR VGND sg13g2_decap_8
XFILLER_82_846 VPWR VGND sg13g2_decap_8
XFILLER_81_323 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_93_194 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q net3323 VGND VPWR i_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[244\] clknet_leaf_56_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y VGND VPWR net1393 net2301 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ net2591 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_50_765 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[8\]_sg13g2_dfrbpq_1_Q net3241 VGND VPWR rsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[8\] clknet_leaf_39_clk sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1065 net697 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\] net649 net2623
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xhold630 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\] VPWR
+ VGND net662 sg13g2_dlygate4sd3_1
Xhold652 data_pdata\[0\] VPWR VGND net684 sg13g2_dlygate4sd3_1
Xhold663 i_snitch.sb_q\[1\] VPWR VGND net695 sg13g2_dlygate4sd3_1
XFILLER_2_817 VPWR VGND sg13g2_decap_8
Xhold641 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_inv_1_A_Y VPWR VGND net673 sg13g2_dlygate4sd3_1
Xfanout2809 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_B net2809 VPWR VGND
+ sg13g2_buf_8
Xhold674 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\] VPWR
+ VGND net706 sg13g2_dlygate4sd3_1
Xhold696 i_snitch.i_snitch_regfile.mem\[127\] VPWR VGND net728 sg13g2_dlygate4sd3_1
Xhold685 i_snitch.i_snitch_regfile.mem\[320\] VPWR VGND net717 sg13g2_dlygate4sd3_1
XFILLER_103_266 VPWR VGND sg13g2_decap_8
XFILLER_77_607 VPWR VGND sg13g2_fill_1
XFILLER_98_990 VPWR VGND sg13g2_decap_8
XFILLER_58_832 VPWR VGND sg13g2_fill_1
XFILLER_58_821 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]
+ net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B net3163 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_2
XFILLER_100_973 VPWR VGND sg13g2_decap_8
XFILLER_94_49 VPWR VGND sg13g2_decap_8
Xhold1341 i_snitch.inst_addr_o\[26\] VPWR VGND net1373 sg13g2_dlygate4sd3_1
Xhold1330 rsp_data_q\[19\] VPWR VGND net1362 sg13g2_dlygate4sd3_1
Xhold1352 rsp_data_q\[21\] VPWR VGND net1384 sg13g2_dlygate4sd3_1
Xhold1363 i_snitch.inst_addr_o\[16\] VPWR VGND net1395 sg13g2_dlygate4sd3_1
Xhold1374 i_snitch.inst_addr_o\[22\] VPWR VGND net1406 sg13g2_dlygate4sd3_1
XFILLER_73_824 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[10\]_sg13g2_nor2_1_A net468 net2733 shift_reg_q\[10\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D
+ net3035 net3147 net2927 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X
+ VPWR VGND sg13g2_and4_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net3032 i_snitch.sb_q\[2\] VPWR VGND sg13g2_nand2b_1
XFILLER_13_412 VPWR VGND sg13g2_decap_4
XFILLER_14_935 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q
+ net3191 VGND VPWR net680 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_25_261 VPWR VGND sg13g2_fill_1
XFILLER_9_405 VPWR VGND sg13g2_fill_2
XFILLER_13_445 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net1010 net2453 net2273 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[369\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net888 net2663 net2883 VPWR VGND sg13g2_a22oi_1
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2321
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q
+ net3247 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_dfrbpq_1_Q net3308 VGND VPWR i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[264\] clknet_leaf_70_clk sg13g2_dfrbpq_1
XFILLER_67_128 VPWR VGND sg13g2_fill_2
XFILLER_49_832 VPWR VGND sg13g2_decap_8
XFILLER_49_821 VPWR VGND sg13g2_fill_1
XFILLER_76_662 VPWR VGND sg13g2_fill_2
XFILLER_0_393 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_76_695 VPWR VGND sg13g2_fill_2
XFILLER_76_684 VPWR VGND sg13g2_fill_1
XFILLER_76_673 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_1_1021 VPWR VGND sg13g2_decap_8
XFILLER_36_559 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y
+ VGND sg13g2_inv_1
XFILLER_91_698 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2334
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ VGND net2707 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
XFILLER_17_784 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2365
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2586 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_949 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y net2519 VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1
+ VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D_sg13g2_nor2_1_Y
+ net75 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D
+ VPWR VGND sg13g2_nor2_1
XFILLER_99_743 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_101_715 VPWR VGND sg13g2_decap_8
XFILLER_87_916 VPWR VGND sg13g2_decap_8
XFILLER_63_1027 VPWR VGND sg13g2_fill_2
XFILLER_101_726 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[23\]_sg13g2_nor2_1_A net511 net2734 shift_reg_q\[23\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_100_247 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR net580 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[39\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_66_161 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2340
+ sg13g2_o21ai_1
XFILLER_10_426 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[65\]
+ net3120 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[284\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2358
+ sg13g2_o21ai_1
XFILLER_6_419 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1 net2527 VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2414
+ sg13g2_o21ai_1
Xfanout3318 net3326 net3318 VPWR VGND sg13g2_buf_8
Xfanout3307 net3311 net3307 VPWR VGND sg13g2_buf_8
XFILLER_2_614 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q
+ net3185 VGND VPWR net607 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
Xfanout3329 net3330 net3329 VPWR VGND sg13g2_buf_8
Xfanout2606 net2607 net2606 VPWR VGND sg13g2_buf_1
Xhold471 shift_reg_q\[8\] VPWR VGND net503 sg13g2_dlygate4sd3_1
Xfanout2617 net2618 net2617 VPWR VGND sg13g2_buf_8
Xhold460 shift_reg_q\[7\] VPWR VGND net492 sg13g2_dlygate4sd3_1
XFILLER_78_938 VPWR VGND sg13g2_decap_8
XFILLER_78_905 VPWR VGND sg13g2_fill_1
Xfanout2628 net2630 net2628 VPWR VGND sg13g2_buf_8
Xhold493 strb_reg_q\[1\] VPWR VGND net525 sg13g2_dlygate4sd3_1
Xhold482 i_snitch.i_snitch_regfile.mem\[33\] VPWR VGND net514 sg13g2_dlygate4sd3_1
Xfanout2639 net2640 net2639 VPWR VGND sg13g2_buf_8
XFILLER_77_437 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2436 net2872 i_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
XFILLER_92_407 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2
+ VPWR VGND sg13g2_nor2_1
XFILLER_86_993 VPWR VGND sg13g2_decap_8
XFILLER_18_504 VPWR VGND sg13g2_decap_8
Xhold1160 i_snitch.i_snitch_regfile.mem\[170\] VPWR VGND net1192 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1369 net2492 net1208 VPWR VGND sg13g2_a22oi_1
Xhold1182 i_snitch.i_snitch_regfile.mem\[445\] VPWR VGND net1214 sg13g2_dlygate4sd3_1
Xhold1193 i_snitch.i_snitch_regfile.mem\[400\] VPWR VGND net1225 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[419\] clknet_leaf_112_clk sg13g2_dfrbpq_1
Xhold1171 i_snitch.i_snitch_regfile.mem\[81\] VPWR VGND net1203 sg13g2_dlygate4sd3_1
XFILLER_45_378 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2858
+ net2656 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2444 VPWR VGND sg13g2_nand2_1
XFILLER_33_507 VPWR VGND sg13g2_fill_2
XFILLER_72_186 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2399
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[208\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net980 net2441 net2263 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]
+ net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_13_242 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_14_798 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q net3215 VGND VPWR i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[103\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ net2627 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xclkload16 clkload16/Y clknet_leaf_16_clk VPWR VGND sg13g2_inv_2
Xclkload27 VPWR clkload27/Y clknet_leaf_21_clk VGND sg13g2_inv_1
Xclkload49 clkload49/Y clknet_leaf_71_clk VPWR VGND sg13g2_inv_2
XFILLER_6_942 VPWR VGND sg13g2_decap_8
Xclkload38 clknet_leaf_103_clk clkload38/X VPWR VGND sg13g2_buf_8
Xi_snitch.wake_up_q\[2\]_sg13g2_nor4_1_D net3 net553 i_snitch.wake_up_q\[0\] net545
+ i_snitch.wake_up_q\[2\]_sg13g2_nor4_1_D_Y VPWR VGND sg13g2_nor4_1
XFILLER_96_757 VPWR VGND sg13g2_decap_8
XFILLER_84_919 VPWR VGND sg13g2_decap_8
XFILLER_0_190 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2748 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_95_278 VPWR VGND sg13g2_fill_2
XFILLER_92_941 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR data_pvalid_sg13g2_dfrbpq_1_Q_D
+ net3052 VGND sg13g2_inv_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B net2626
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_64_665 VPWR VGND sg13g2_fill_2
Xdata_pdata\[7\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B net3153 data_pdata\[7\]_sg13g2_mux2_1_A0_X
+ data_pdata\[7\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D
+ net915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_52_838 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0 net3130 i_snitch.i_snitch_regfile.mem\[142\]
+ i_snitch.i_snitch_regfile.mem\[174\] i_snitch.i_snitch_regfile.mem\[206\] i_snitch.i_snitch_regfile.mem\[238\]
+ net3109 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2860
+ net2673 VPWR VGND sg13g2_nand2_1
XFILLER_81_0 VPWR VGND sg13g2_decap_8
XFILLER_20_735 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2594 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1_sg13g2_o21ai_1_Y
+ net2549 VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1
+ VGND net2715 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
XFILLER_106_829 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A
+ net36 net2509 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_99_562 VPWR VGND sg13g2_decap_4
XFILLER_99_540 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[439\] clknet_leaf_67_clk sg13g2_dfrbpq_1
XFILLER_101_545 VPWR VGND sg13g2_fill_1
XFILLER_101_534 VPWR VGND sg13g2_decap_8
XFILLER_87_768 VPWR VGND sg13g2_fill_1
XFILLER_101_589 VPWR VGND sg13g2_fill_1
XFILLER_101_578 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ net2696 VPWR VGND sg13g2_inv_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]
+ net3171 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_55_610 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1133 net869 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[123\] clknet_leaf_112_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2891 net2906 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_83_963 VPWR VGND sg13g2_decap_8
XFILLER_82_451 VPWR VGND sg13g2_fill_1
XFILLER_70_602 VPWR VGND sg13g2_fill_2
XFILLER_55_676 VPWR VGND sg13g2_fill_1
XFILLER_55_654 VPWR VGND sg13g2_fill_2
XFILLER_91_28 VPWR VGND sg13g2_decap_4
XFILLER_43_849 VPWR VGND sg13g2_decap_4
XFILLER_43_838 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0 net3118 i_snitch.i_snitch_regfile.mem\[261\]
+ i_snitch.i_snitch_regfile.mem\[293\] i_snitch.i_snitch_regfile.mem\[325\] i_snitch.i_snitch_regfile.mem\[357\]
+ net3102 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_36_890 VPWR VGND sg13g2_fill_1
Xi_req_arb.data_i\[42\]_sg13g2_dfrbpq_1_Q net3260 VGND VPWR i_snitch.pc_d\[7\] i_req_arb.data_i\[42\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_23_573 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2881
+ net2693 VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[22\]_sg13g2_dfrbpq_1_Q net3200 VGND VPWR net542 shift_reg_q\[22\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_10_289 VPWR VGND sg13g2_fill_2
Xfanout3104 net3105 net3104 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B net2816
+ i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_105_840 VPWR VGND sg13g2_decap_8
Xfanout3137 net3139 net3137 VPWR VGND sg13g2_buf_8
XFILLER_3_934 VPWR VGND sg13g2_decap_8
Xfanout3115 net3118 net3115 VPWR VGND sg13g2_buf_8
Xfanout3126 net3128 net3126 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[81\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[81\]
+ i_snitch.i_snitch_regfile.mem\[113\] net3130 i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_104_350 VPWR VGND sg13g2_decap_8
Xfanout3148 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1_X
+ net3148 VPWR VGND sg13g2_buf_8
Xfanout2414 i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ net2414 VPWR VGND sg13g2_buf_8
Xfanout2425 net2427 net2425 VPWR VGND sg13g2_buf_8
Xfanout3159 net3160 net3159 VPWR VGND sg13g2_buf_2
Xfanout2403 net2406 net2403 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2629 net2761 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2742
+ net2675 VPWR VGND sg13g2_nand2_1
Xfanout2469 net2471 net2469 VPWR VGND sg13g2_buf_8
Xfanout2458 net2459 net2458 VPWR VGND sg13g2_buf_8
Xfanout2436 net2438 net2436 VPWR VGND sg13g2_buf_8
Xfanout2447 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2447 VPWR
+ VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2490 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor2_1_B
+ net3107 net2953 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_A2 VPWR VGND
+ sg13g2_nor2_2
XFILLER_93_716 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B
+ net2566 sg13g2_a21oi_1
Xi_req_arb.data_i\[37\]_sg13g2_inv_1_A i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_A i_req_arb.data_i\[37\]
+ VPWR VGND sg13g2_inv_2
XFILLER_105_91 VPWR VGND sg13g2_decap_8
XFILLER_58_481 VPWR VGND sg13g2_fill_1
XFILLER_19_846 VPWR VGND sg13g2_decap_4
XFILLER_46_698 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2462
+ net2283 net2694 net2742 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2592 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2698 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ net2540 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[459\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[248\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[248\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net899 net2666 net2875 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_53_4 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C
+ VPWR i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2
+ VGND net2565 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ net2526 i_snitch.inst_addr_o\[23\] sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q net3299 VGND VPWR i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[143\] clknet_leaf_63_clk sg13g2_dfrbpq_1
Xfanout2981 net2984 net2981 VPWR VGND sg13g2_buf_1
Xfanout2970 net2972 net2970 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y
+ net53 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ sg13g2_a21oi_2
XFILLER_56_418 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_mux4_1_X
+ net3122 i_snitch.sb_q\[4\] i_snitch.sb_q\[5\] i_snitch.sb_q\[6\] i_snitch.sb_q\[7\]
+ net3104 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux4_1
Xfanout2992 net2994 net2992 VPWR VGND sg13g2_buf_8
XFILLER_84_749 VPWR VGND sg13g2_decap_4
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_nor2_1_A net692 net2488 i_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_92_771 VPWR VGND sg13g2_fill_1
XFILLER_91_281 VPWR VGND sg13g2_fill_2
XFILLER_64_473 VPWR VGND sg13g2_fill_1
XFILLER_101_49 VPWR VGND sg13g2_decap_8
XFILLER_80_966 VPWR VGND sg13g2_decap_8
XFILLER_52_657 VPWR VGND sg13g2_fill_2
XFILLER_52_646 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2467
+ net2514 net2902 net3040 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y
+ net432 VGND sg13g2_inv_1
XFILLER_32_381 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[471\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[471\] net2952 VPWR VGND sg13g2_nand2_1
XFILLER_20_598 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y net2637
+ sg13g2_a21oi_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_mux4_1_X
+ net3007 i_snitch.sb_q\[12\] i_snitch.sb_q\[13\] i_snitch.sb_q\[14\] i_snitch.sb_q\[15\]
+ net2980 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_mux4_1
XFILLER_3_219 VPWR VGND sg13g2_fill_2
XFILLER_105_147 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[6\]_sg13g2_nor2b_1_A i_snitch.gpr_waddr\[6\] i_snitch.gpr_waddr\[7\]
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B VPWR
+ VGND sg13g2_nor2b_2
XFILLER_102_821 VPWR VGND sg13g2_decap_8
XFILLER_0_926 VPWR VGND sg13g2_decap_8
XFILLER_102_898 VPWR VGND sg13g2_decap_8
XFILLER_101_364 VPWR VGND sg13g2_decap_8
XFILLER_87_576 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_fill_1
XFILLER_74_237 VPWR VGND sg13g2_fill_2
XFILLER_28_610 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2879
+ i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand3_1_C
+ net119 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_76_1004 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y
+ net2932 net3096 VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[479\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_83_793 VPWR VGND sg13g2_decap_8
XFILLER_70_421 VPWR VGND sg13g2_fill_2
XFILLER_43_613 VPWR VGND sg13g2_fill_1
XFILLER_27_164 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[268\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2326 net811 net2691 net2894 VPWR VGND sg13g2_a22oi_1
XFILLER_15_348 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0 net3119 i_snitch.i_snitch_regfile.mem\[149\]
+ i_snitch.i_snitch_regfile.mem\[181\] i_snitch.i_snitch_regfile.mem\[213\] i_snitch.i_snitch_regfile.mem\[245\]
+ net3101 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xclkbuf_leaf_116_clk clknet_5_5__leaf_clk clknet_leaf_116_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[163\] clknet_leaf_108_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2713 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nor2b_1
XFILLER_7_525 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0_1 i_snitch.i_snitch_regfile.mem\[193\]
+ i_snitch.i_snitch_regfile.mem\[225\] net3133 i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_98_808 VPWR VGND sg13g2_decap_8
Xi_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y VGND
+ VPWR net553 i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C net545 sg13g2_a21oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xnor2_1
XFILLER_83_1019 VPWR VGND sg13g2_decap_8
Xfanout2244 net2245 net2244 VPWR VGND sg13g2_buf_8
Xfanout2277 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_Y
+ net2277 VPWR VGND sg13g2_buf_8
Xfanout2266 net2267 net2266 VPWR VGND sg13g2_buf_8
Xfanout2255 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2255 VPWR VGND sg13g2_buf_8
XFILLER_93_502 VPWR VGND sg13g2_decap_8
Xfanout2299 net2300 net2299 VPWR VGND sg13g2_buf_8
Xfanout2288 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2288 VPWR VGND sg13g2_buf_8
XFILLER_74_760 VPWR VGND sg13g2_decap_8
XFILLER_20_1025 VPWR VGND sg13g2_decap_4
XFILLER_18_197 VPWR VGND sg13g2_decap_4
XFILLER_22_819 VPWR VGND sg13g2_decap_4
XFILLER_15_893 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_107_clk clknet_5_7__leaf_clk clknet_leaf_107_clk VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y
+ net445 VGND sg13g2_inv_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A
+ net2707 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y
+ net2925 net2926 net3033 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A
+ VPWR VGND net2922 sg13g2_nand4_1
XFILLER_103_629 VPWR VGND sg13g2_fill_1
XFILLER_103_618 VPWR VGND sg13g2_decap_4
XFILLER_88_318 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[499\] clknet_leaf_116_clk sg13g2_dfrbpq_1
XFILLER_97_852 VPWR VGND sg13g2_decap_8
XFILLER_69_554 VPWR VGND sg13g2_fill_2
XFILLER_69_532 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2729 shift_reg_q\[21\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[17\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[17\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[278\] net3029 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[288\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2904 net2778 net2316 net1254 VPWR VGND sg13g2_a22oi_1
XFILLER_5_1019 VPWR VGND sg13g2_decap_8
XFILLER_84_546 VPWR VGND sg13g2_decap_4
XFILLER_57_738 VPWR VGND sg13g2_fill_1
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_72_708 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C
+ net2429 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_37_440 VPWR VGND sg13g2_fill_1
XFILLER_37_451 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[183\] clknet_leaf_57_clk sg13g2_dfrbpq_1
XFILLER_65_782 VPWR VGND sg13g2_fill_2
XFILLER_65_771 VPWR VGND sg13g2_decap_8
XFILLER_53_922 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[387\] VGND sg13g2_inv_1
XFILLER_25_624 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B
+ net2701 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_33_690 VPWR VGND sg13g2_fill_2
XFILLER_20_351 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0 net3121 i_snitch.i_snitch_regfile.mem\[387\]
+ i_snitch.i_snitch_regfile.mem\[419\] i_snitch.i_snitch_regfile.mem\[451\] i_snitch.i_snitch_regfile.mem\[483\]
+ net3101 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_106_434 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[318\] clknet_leaf_94_clk sg13g2_dfrbpq_1
XFILLER_97_49 VPWR VGND sg13g2_decap_8
XFILLER_0_723 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[107\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net817 net2680 net2871 VPWR VGND sg13g2_a22oi_1
XFILLER_102_662 VPWR VGND sg13g2_fill_1
XFILLER_88_896 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[1\]_sg13g2_dfrbpq_1_Q net3185 VGND VPWR net526 strb_reg_q\[1\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
XFILLER_102_695 VPWR VGND sg13g2_decap_8
XFILLER_101_161 VPWR VGND sg13g2_decap_8
XFILLER_75_546 VPWR VGND sg13g2_decap_4
Xdata_pdata\[15\]_sg13g2_mux2_1_A1 rsp_data_q\[15\] net966 net3052 data_pdata\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_75_579 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_55_270 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2475 net2466 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2
+ VGND VPWR net2711 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_B
+ net2612 sg13g2_a21oi_1
XFILLER_90_549 VPWR VGND sg13g2_fill_1
XFILLER_46_97 VPWR VGND sg13g2_decap_4
XFILLER_102_70 VPWR VGND sg13g2_decap_8
XFILLER_15_167 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
XFILLER_50_1018 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_fill_1
XFILLER_8_845 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_4
XFILLER_7_25 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y
+ net441 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1
+ VPWR VGND sg13g2_nor3_1
XFILLER_106_990 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_o21ai_1_A1 net2970 VPWR i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[370\] net2805 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_93_321 VPWR VGND sg13g2_fill_1
XFILLER_78_395 VPWR VGND sg13g2_decap_8
XFILLER_93_354 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[51\] clknet_leaf_113_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VGND i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ sg13g2_o21ai_1
XFILLER_35_944 VPWR VGND sg13g2_fill_2
XFILLER_62_785 VPWR VGND sg13g2_fill_1
XFILLER_62_763 VPWR VGND sg13g2_fill_2
XFILLER_21_126 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[338\] clknet_leaf_91_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[127\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2410 net728 net2646 net2869 VPWR VGND sg13g2_a22oi_1
Xhold801 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] VPWR
+ VGND net833 sg13g2_dlygate4sd3_1
Xhold812 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\] VPWR
+ VGND net844 sg13g2_dlygate4sd3_1
Xhold834 i_snitch.i_snitch_regfile.mem\[180\] VPWR VGND net866 sg13g2_dlygate4sd3_1
Xhold823 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net855 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_o21ai_1_A1 net3023 VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[47\] net2994 sg13g2_o21ai_1
Xhold845 i_snitch.i_snitch_regfile.mem\[85\] VPWR VGND net877 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1 net3117 i_snitch.i_snitch_regfile.mem\[130\]
+ i_snitch.i_snitch_regfile.mem\[162\] i_snitch.i_snitch_regfile.mem\[194\] i_snitch.i_snitch_regfile.mem\[226\]
+ net3099 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_104_949 VPWR VGND sg13g2_decap_8
XFILLER_103_415 VPWR VGND sg13g2_fill_1
Xhold867 i_snitch.i_snitch_regfile.mem\[248\] VPWR VGND net899 sg13g2_dlygate4sd3_1
Xhold878 i_snitch.i_snitch_regfile.mem\[160\] VPWR VGND net910 sg13g2_dlygate4sd3_1
Xhold856 i_snitch.i_snitch_regfile.mem\[369\] VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold889 i_snitch.i_snitch_regfile.mem\[254\] VPWR VGND net921 sg13g2_dlygate4sd3_1
Xshift_reg_q\[26\]_sg13g2_a22oi_1_A1 shift_reg_q\[26\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[32\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[26\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\] clknet_leaf_47_clk
+ sg13g2_dfrbpq_1
XFILLER_85_899 VPWR VGND sg13g2_decap_8
XFILLER_38_760 VPWR VGND sg13g2_decap_4
XFILLER_37_270 VPWR VGND sg13g2_decap_8
XFILLER_52_240 VPWR VGND sg13g2_fill_1
XFILLER_16_45 VPWR VGND sg13g2_fill_2
XFILLER_40_402 VPWR VGND sg13g2_decap_8
XFILLER_52_273 VPWR VGND sg13g2_decap_8
XFILLER_40_435 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]
+ net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X
+ VPWR VGND sg13g2_or4_1
XFILLER_32_77 VPWR VGND sg13g2_fill_1
XFILLER_10_1013 VPWR VGND sg13g2_decap_8
XFILLER_106_231 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C i_snitch.inst_addr_o\[17\]
+ net2306 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[71\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2542 VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VGND net2750 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C
+ net2710 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X
+ VPWR VGND sg13g2_or4_1
XFILLER_76_811 VPWR VGND sg13g2_fill_2
XFILLER_102_481 VPWR VGND sg13g2_fill_2
XFILLER_102_470 VPWR VGND sg13g2_decap_8
XFILLER_88_693 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ sg13g2_a21oi_1
XFILLER_48_513 VPWR VGND sg13g2_decap_8
XFILLER_0_597 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_48_579 VPWR VGND sg13g2_decap_4
XFILLER_36_719 VPWR VGND sg13g2_fill_2
XFILLER_17_900 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[358\] clknet_leaf_77_clk sg13g2_dfrbpq_1
XFILLER_90_357 VPWR VGND sg13g2_decap_8
XFILLER_17_933 VPWR VGND sg13g2_decap_8
XFILLER_90_368 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_44_785 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net1033 net2445 net2270 VPWR VGND sg13g2_a22oi_1
XFILLER_32_947 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1 net3122 i_snitch.i_snitch_regfile.mem\[132\]
+ i_snitch.i_snitch_regfile.mem\[164\] i_snitch.i_snitch_regfile.mem\[196\] i_snitch.i_snitch_regfile.mem\[228\]
+ net3104 i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_671 VPWR VGND sg13g2_decap_8
XFILLER_89_1014 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A
+ net3144 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_98_70 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D
+ net2744 net2928 sg13g2_a21oi_2
XFILLER_99_958 VPWR VGND sg13g2_decap_8
XFILLER_67_800 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_94_652 VPWR VGND sg13g2_decap_4
Xi_snitch.inst_addr_o\[18\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[18\]
+ i_snitch.inst_addr_o\[18\] clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_67_855 VPWR VGND sg13g2_decap_4
XFILLER_94_674 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1126 net1063 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_26_207 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B_sg13g2_and2_1_X net1391 net3172 i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B
+ VPWR VGND sg13g2_and2_1
XFILLER_22_479 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[91\] clknet_leaf_112_clk sg13g2_dfrbpq_1
XFILLER_30_490 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q
+ net3238 VGND VPWR net773 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2400
+ sg13g2_o21ai_1
Xhold620 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net652 sg13g2_dlygate4sd3_1
XFILLER_104_702 VPWR VGND sg13g2_fill_2
Xhold653 data_pdata\[0\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net685 sg13g2_dlygate4sd3_1
Xhold631 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net663 sg13g2_dlygate4sd3_1
Xhold642 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y VPWR VGND net674 sg13g2_dlygate4sd3_1
Xhold664 i_snitch.inst_addr_o\[31\] VPWR VGND net696 sg13g2_dlygate4sd3_1
Xhold686 i_snitch.i_snitch_regfile.mem\[212\] VPWR VGND net718 sg13g2_dlygate4sd3_1
Xhold675 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net707 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[378\] clknet_leaf_115_clk sg13g2_dfrbpq_1
Xhold697 data_pdata\[17\] VPWR VGND net729 sg13g2_dlygate4sd3_1
XFILLER_103_245 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[167\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2442 net2284 net2342 net1163 VPWR VGND sg13g2_a22oi_1
XFILLER_100_952 VPWR VGND sg13g2_decap_8
XFILLER_94_28 VPWR VGND sg13g2_decap_8
Xhold1331 i_snitch.inst_addr_o\[14\] VPWR VGND net1363 sg13g2_dlygate4sd3_1
Xhold1342 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] VPWR
+ VGND net1374 sg13g2_dlygate4sd3_1
Xhold1320 i_snitch.i_snitch_regfile.mem\[55\] VPWR VGND net1352 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_96_clk clknet_5_17__leaf_clk clknet_leaf_96_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1 net3013 i_snitch.i_snitch_regfile.mem\[134\]
+ i_snitch.i_snitch_regfile.mem\[166\] i_snitch.i_snitch_regfile.mem\[198\] i_snitch.i_snitch_regfile.mem\[230\]
+ net2986 i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
XFILLER_85_674 VPWR VGND sg13g2_fill_1
Xhold1353 i_snitch.inst_addr_o\[11\] VPWR VGND net1385 sg13g2_dlygate4sd3_1
Xhold1364 i_snitch.inst_addr_o\[15\] VPWR VGND net1396 sg13g2_dlygate4sd3_1
Xhold1375 i_snitch.i_snitch_lsu.handshake_pending_q VPWR VGND net1407 sg13g2_dlygate4sd3_1
XFILLER_58_899 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B sg13g2_o21ai_1
XFILLER_72_335 VPWR VGND sg13g2_decap_4
XFILLER_27_77 VPWR VGND sg13g2_fill_2
XFILLER_26_752 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2445 net2887 i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
XFILLER_26_785 VPWR VGND sg13g2_fill_1
XFILLER_26_796 VPWR VGND sg13g2_fill_2
XFILLER_41_711 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[4\]_sg13g2_nor2_1_A net465 net2736 shift_reg_q\[4\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2480 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[122\]
+ net2998 i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_40_276 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_20_clk clknet_5_12__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_4_133 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2281
+ sg13g2_o21ai_1
XFILLER_68_40 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_67_107 VPWR VGND sg13g2_fill_2
XFILLER_0_372 VPWR VGND sg13g2_decap_8
XFILLER_1_895 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_87_clk clknet_5_21__leaf_clk clknet_leaf_87_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D_sg13g2_or2_1_X
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ net3087 sg13g2_or2_1
XFILLER_63_302 VPWR VGND sg13g2_fill_2
XFILLER_49_888 VPWR VGND sg13g2_decap_8
XFILLER_48_387 VPWR VGND sg13g2_fill_2
XFILLER_1_1000 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1293 net3065 rsp_data_q\[25\] VPWR VGND sg13g2_a22oi_1
XFILLER_64_858 VPWR VGND sg13g2_decap_4
XFILLER_48_398 VPWR VGND sg13g2_decap_8
XFILLER_91_688 VPWR VGND sg13g2_fill_1
XFILLER_91_677 VPWR VGND sg13g2_fill_2
XFILLER_91_666 VPWR VGND sg13g2_fill_2
XFILLER_51_519 VPWR VGND sg13g2_fill_1
XFILLER_90_198 VPWR VGND sg13g2_fill_2
XFILLER_31_232 VPWR VGND sg13g2_decap_4
XFILLER_83_4 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q
+ net3250 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
XFILLER_20_939 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_11_clk clknet_5_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[398\] clknet_leaf_78_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_or3_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_B
+ VPWR VGND sg13g2_or3_1
Xi_snitch.i_snitch_regfile.mem\[187\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2442 net2252 net2342 net1278 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2696 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_mux2_1_A1
+ net991 net563 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1 net3008 i_snitch.i_snitch_regfile.mem\[136\]
+ i_snitch.i_snitch_regfile.mem\[168\] i_snitch.i_snitch_regfile.mem\[200\] i_snitch.i_snitch_regfile.mem\[232\]
+ net2982 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2377
+ sg13g2_o21ai_1
XFILLER_100_226 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_mux2_1_A0_X net3101 net2824 i_snitch.i_snitch_regfile.mem\[35\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_78_clk clknet_5_22__leaf_clk clknet_leaf_78_clk VPWR VGND sg13g2_buf_8
XFILLER_39_332 VPWR VGND sg13g2_fill_2
XFILLER_104_49 VPWR VGND sg13g2_decap_8
XFILLER_95_994 VPWR VGND sg13g2_decap_8
XFILLER_39_354 VPWR VGND sg13g2_fill_1
XFILLER_94_493 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2385
+ sg13g2_o21ai_1
XFILLER_55_858 VPWR VGND sg13g2_fill_2
XFILLER_70_806 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1
+ net2547 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B
+ sg13g2_a221oi_1
XFILLER_23_744 VPWR VGND sg13g2_fill_1
XFILLER_10_405 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[217\] clknet_leaf_116_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_23_788 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[36\]
+ net3008 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1_Y net2980 sg13g2_a21oi_1
Xfanout3319 net3325 net3319 VPWR VGND sg13g2_buf_8
Xfanout3308 net3311 net3308 VPWR VGND sg13g2_buf_8
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y i_snitch.gpr_waddr\[6\]
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.gpr_waddr\[7\]
+ i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand3_1
Xfanout2607 net65 net2607 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net123 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y
+ net553 net545 i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
Xhold472 shift_reg_q\[8\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold450 shift_reg_q\[17\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net482 sg13g2_dlygate4sd3_1
Xfanout2618 net2620 net2618 VPWR VGND sg13g2_buf_8
Xhold461 shift_reg_q\[7\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net493 sg13g2_dlygate4sd3_1
Xfanout2629 net2630 net2629 VPWR VGND sg13g2_buf_8
XFILLER_1_147 VPWR VGND sg13g2_decap_4
Xhold494 strb_reg_q\[1\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net526 sg13g2_dlygate4sd3_1
Xshift_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2730 shift_reg_q\[9\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[5\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold483 shift_reg_q\[25\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2364
+ sg13g2_o21ai_1
XFILLER_49_129 VPWR VGND sg13g2_decap_4
XFILLER_93_909 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_69_clk clknet_5_27__leaf_clk clknet_leaf_69_clk VPWR VGND sg13g2_buf_8
XFILLER_86_972 VPWR VGND sg13g2_decap_8
XFILLER_85_460 VPWR VGND sg13g2_fill_2
Xhold1150 i_snitch.i_snitch_regfile.mem\[311\] VPWR VGND net1182 sg13g2_dlygate4sd3_1
Xhold1194 rsp_data_q\[18\] VPWR VGND net1226 sg13g2_dlygate4sd3_1
Xhold1161 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] VPWR
+ VGND net1193 sg13g2_dlygate4sd3_1
XFILLER_45_335 VPWR VGND sg13g2_decap_4
XFILLER_45_313 VPWR VGND sg13g2_fill_2
Xhold1183 i_snitch.i_snitch_regfile.mem\[186\] VPWR VGND net1215 sg13g2_dlygate4sd3_1
Xhold1172 i_snitch.i_snitch_regfile.mem\[117\] VPWR VGND net1204 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2596 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_73_677 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2496 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_33_519 VPWR VGND sg13g2_fill_2
XFILLER_72_176 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2392
+ sg13g2_o21ai_1
XFILLER_14_733 VPWR VGND sg13g2_fill_1
XFILLER_13_221 VPWR VGND sg13g2_decap_4
XFILLER_14_744 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1 net3014 i_snitch.i_snitch_regfile.mem\[138\]
+ i_snitch.i_snitch_regfile.mem\[170\] i_snitch.i_snitch_regfile.mem\[202\] i_snitch.i_snitch_regfile.mem\[234\]
+ net2986 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_6_921 VPWR VGND sg13g2_decap_8
Xclkload17 clknet_leaf_107_clk clkload17/X VPWR VGND sg13g2_buf_8
Xclkload28 clknet_leaf_22_clk clkload28/Y VPWR VGND sg13g2_inv_4
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_mux2_1_A0_X net3111 net2829 i_snitch.i_snitch_regfile.mem\[55\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net1352 net2648 net2769 VPWR VGND sg13g2_a22oi_1
Xclkload39 clkload39/Y clknet_leaf_92_clk VPWR VGND sg13g2_inv_2
XFILLER_86_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_998 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1 net3117 i_snitch.i_snitch_regfile.mem\[386\]
+ i_snitch.i_snitch_regfile.mem\[418\] i_snitch.i_snitch_regfile.mem\[450\] i_snitch.i_snitch_regfile.mem\[482\]
+ net3102 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_96_714 VPWR VGND sg13g2_fill_1
XFILLER_1_692 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_92_920 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[56\]
+ net2828 i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a21oi_1_A1_Y net2823 sg13g2_a21oi_1
Xclkbuf_leaf_0_clk clknet_5_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net514 net2359 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[237\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_37_847 VPWR VGND sg13g2_decap_4
XFILLER_91_441 VPWR VGND sg13g2_decap_4
XFILLER_92_997 VPWR VGND sg13g2_decap_8
XFILLER_45_880 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A_sg13g2_or2_1_X
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2566 sg13g2_or2_1
XFILLER_60_861 VPWR VGND sg13g2_fill_1
XFILLER_20_714 VPWR VGND sg13g2_decap_8
XFILLER_32_563 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2450 VPWR VGND sg13g2_nand2_1
XFILLER_106_808 VPWR VGND sg13g2_decap_8
XFILLER_105_329 VPWR VGND sg13g2_decap_8
XFILLER_99_552 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y net2724
+ net2955 VPWR VGND sg13g2_a22oi_1
XFILLER_83_942 VPWR VGND sg13g2_decap_8
XFILLER_67_493 VPWR VGND sg13g2_fill_2
XFILLER_28_836 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 VGND sg13g2_inv_1
XFILLER_27_357 VPWR VGND sg13g2_fill_1
XFILLER_55_699 VPWR VGND sg13g2_decap_4
XFILLER_42_327 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[75\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net934 net2679 net2787 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\] net625 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2781
+ net2650 VPWR VGND sg13g2_nand2_1
XFILLER_3_913 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2415 sg13g2_a21oi_1
Xfanout3105 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_X
+ net3105 VPWR VGND sg13g2_buf_8
Xfanout3138 net3139 net3138 VPWR VGND sg13g2_buf_8
Xfanout3116 net3118 net3116 VPWR VGND sg13g2_buf_8
Xfanout3127 net3128 net3127 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[257\] clknet_leaf_103_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0
+ sg13g2_a21oi_1
XFILLER_78_703 VPWR VGND sg13g2_fill_2
Xfanout2426 net2427 net2426 VPWR VGND sg13g2_buf_8
XFILLER_46_1023 VPWR VGND sg13g2_decap_4
Xfanout2415 net2416 net2415 VPWR VGND sg13g2_buf_2
Xfanout3149 net3150 net3149 VPWR VGND sg13g2_buf_8
Xfanout2404 net2405 net2404 VPWR VGND sg13g2_buf_1
XFILLER_105_896 VPWR VGND sg13g2_decap_8
Xfanout2448 net2449 net2448 VPWR VGND sg13g2_buf_8
Xfanout2437 net2438 net2437 VPWR VGND sg13g2_buf_8
Xfanout2459 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2459 VPWR
+ VGND sg13g2_buf_8
XFILLER_78_758 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2446 VPWR VGND sg13g2_nand2_1
XFILLER_105_70 VPWR VGND sg13g2_decap_8
XFILLER_100_590 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2483 VPWR VGND sg13g2_a22oi_1
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_836 VPWR VGND sg13g2_fill_1
XFILLER_19_858 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2
+ net2569 VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ VGND net33 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_45_154 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2334
+ sg13g2_o21ai_1
XFILLER_34_828 VPWR VGND sg13g2_fill_1
XFILLER_14_552 VPWR VGND sg13g2_fill_1
XFILLER_42_872 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2586 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2873
+ net2669 VPWR VGND sg13g2_nand2_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y
+ net2848 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2 VPWR VGND
+ sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2724 i_snitch.inst_addr_o\[13\] sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2828
+ sg13g2_a221oi_1
XFILLER_46_4 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1
+ net2506 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_96_500 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2363
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2798
+ net2653 VPWR VGND sg13g2_nand2_1
XFILLER_96_533 VPWR VGND sg13g2_fill_1
Xfanout2960 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2960 VPWR VGND sg13g2_buf_8
Xfanout2982 net2984 net2982 VPWR VGND sg13g2_buf_8
Xfanout2971 net2972 net2971 VPWR VGND sg13g2_buf_8
XFILLER_84_728 VPWR VGND sg13g2_decap_8
XFILLER_84_717 VPWR VGND sg13g2_decap_8
Xfanout2993 net2994 net2993 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[95\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2354 net731 net2646 net2785 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2747 net2556 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_77_780 VPWR VGND sg13g2_fill_1
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_49_482 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3040
+ net2675 VPWR VGND sg13g2_nand2_1
XFILLER_92_750 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2706 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_80_945 VPWR VGND sg13g2_decap_8
XFILLER_64_485 VPWR VGND sg13g2_fill_2
XFILLER_36_165 VPWR VGND sg13g2_decap_4
XFILLER_101_28 VPWR VGND sg13g2_decap_8
XFILLER_51_135 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ net89 sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y net2753
+ net3080 VPWR VGND sg13g2_a22oi_1
XFILLER_51_168 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q net3264 VGND VPWR i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[277\] clknet_leaf_113_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2854
+ net2659 VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q
+ net3235 VGND VPWR net1127 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_106_638 VPWR VGND sg13g2_fill_2
XFILLER_105_126 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2603 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_0_905 VPWR VGND sg13g2_decap_8
XFILLER_102_800 VPWR VGND sg13g2_decap_8
XFILLER_87_511 VPWR VGND sg13g2_decap_8
XFILLER_87_500 VPWR VGND sg13g2_fill_2
XFILLER_86_29 VPWR VGND sg13g2_decap_8
XFILLER_99_393 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2
+ net2518 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_a21o_1
XFILLER_102_877 VPWR VGND sg13g2_decap_8
XFILLER_101_343 VPWR VGND sg13g2_decap_8
XFILLER_75_706 VPWR VGND sg13g2_decap_8
XFILLER_59_268 VPWR VGND sg13g2_decap_4
XFILLER_74_216 VPWR VGND sg13g2_fill_1
XFILLER_19_67 VPWR VGND sg13g2_decap_4
XFILLER_56_953 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[5\] net998 net2916 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_43_603 VPWR VGND sg13g2_decap_4
XFILLER_15_316 VPWR VGND sg13g2_decap_4
XFILLER_16_839 VPWR VGND sg13g2_fill_1
XFILLER_42_102 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2705 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y
+ VPWR VGND i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D
+ sg13g2_nand4_1
XFILLER_82_282 VPWR VGND sg13g2_fill_2
XFILLER_24_861 VPWR VGND sg13g2_fill_1
XFILLER_42_157 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1362 net2492 net1207 VPWR VGND sg13g2_a22oi_1
XFILLER_23_360 VPWR VGND sg13g2_fill_1
XFILLER_11_555 VPWR VGND sg13g2_fill_2
XFILLER_11_588 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2473
+ net2513 net2901 net2796 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_q\[13\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.sb_d\[13\] i_snitch.sb_q\[13\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_2
Xdata_pdata\[11\]_sg13g2_nand2b_1_B data_pdata\[11\]_sg13g2_nand2b_1_B_Y data_pdata\[11\]
+ net3158 VPWR VGND sg13g2_nand2b_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_3_765 VPWR VGND sg13g2_decap_8
Xfanout2256 net2257 net2256 VPWR VGND sg13g2_buf_8
Xfanout2267 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y
+ net2267 VPWR VGND sg13g2_buf_8
Xfanout2245 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2245 VPWR VGND sg13g2_buf_8
XFILLER_76_40 VPWR VGND sg13g2_fill_1
Xfanout2278 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y
+ net2278 VPWR VGND sg13g2_buf_8
Xfanout2289 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2289 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR
+ VGND net2831 net2638 i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1_Y net2954
+ i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ sg13g2_a221oi_1
XFILLER_65_227 VPWR VGND sg13g2_fill_2
XFILLER_47_953 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[297\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_19_699 VPWR VGND sg13g2_fill_1
XFILLER_61_433 VPWR VGND sg13g2_fill_1
Xdata_pdata\[10\]_sg13g2_dfrbpq_1_Q net3196 VGND VPWR net825 data_pdata\[10\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2606 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VGND net2586 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_33_179 VPWR VGND sg13g2_fill_2
XFILLER_30_842 VPWR VGND sg13g2_fill_1
Xdata_pvalid_sg13g2_nor2_1_A net423 data_pvalid_sg13g2_nor2_1_A_B data_pvalid_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_570 VPWR VGND sg13g2_fill_2
XFILLER_97_831 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0 net3116 i_snitch.i_snitch_regfile.mem\[153\]
+ i_snitch.i_snitch_regfile.mem\[185\] i_snitch.i_snitch_regfile.mem\[217\] i_snitch.i_snitch_regfile.mem\[249\]
+ net3098 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C i_snitch.i_snitch_lsu.metadata_q\[1\]
+ data_pdata\[18\]_sg13g2_mux2_1_A0_X data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y
+ VPWR VGND net3150 sg13g2_nand3b_1
XFILLER_37_0 VPWR VGND sg13g2_fill_1
Xfanout2790 net2793 net2790 VPWR VGND sg13g2_buf_8
XFILLER_96_396 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[116\] clknet_leaf_60_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_nor2b_1_B_N net3115 i_snitch.i_snitch_regfile.mem\[347\]
+ i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_nor2b_1_B_N_Y VPWR VGND sg13g2_nor2b_1
XFILLER_53_901 VPWR VGND sg13g2_decap_4
XFILLER_2_81 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2742
+ net2667 VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3062 net1345 net3065 net1271 VPWR VGND sg13g2_a22oi_1
XFILLER_52_444 VPWR VGND sg13g2_fill_1
XFILLER_52_422 VPWR VGND sg13g2_decap_4
XFILLER_24_113 VPWR VGND sg13g2_fill_1
Xdata_pdata\[31\]_sg13g2_nand2b_1_B data_pdata\[31\]_sg13g2_nand2b_1_B_Y data_pdata\[31\]
+ net3159 VPWR VGND sg13g2_nand2b_1
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[15\]_sg13g2_dfrbpq_1_Q net3197 VGND VPWR net462 shift_reg_q\[15\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_106_413 VPWR VGND sg13g2_decap_8
XFILLER_21_68 VPWR VGND sg13g2_fill_2
XFILLER_97_28 VPWR VGND sg13g2_decap_8
XFILLER_0_702 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2768
+ net2650 VPWR VGND sg13g2_nand2_1
XFILLER_102_674 VPWR VGND sg13g2_fill_1
XFILLER_101_140 VPWR VGND sg13g2_decap_8
XFILLER_88_875 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
Xdata_pdata\[30\]_sg13g2_dfrbpq_1_Q net3204 VGND VPWR net1055 data_pdata\[30\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2467 net2246 net2389 net1129 VPWR VGND sg13g2_a22oi_1
XFILLER_0_779 VPWR VGND sg13g2_decap_8
XFILLER_47_216 VPWR VGND sg13g2_decap_4
XFILLER_47_249 VPWR VGND sg13g2_fill_1
XFILLER_29_942 VPWR VGND sg13g2_fill_1
XFILLER_29_975 VPWR VGND sg13g2_fill_2
XFILLER_90_517 VPWR VGND sg13g2_decap_4
XFILLER_44_901 VPWR VGND sg13g2_fill_2
XFILLER_83_580 VPWR VGND sg13g2_decap_8
XFILLER_43_444 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2897 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ VGND net75 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
XFILLER_70_230 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_820 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[413\]
+ net3028 i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_a21oi_1_A1_Y net2985 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.inst_addr_o\[23\] net2722 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y
+ sg13g2_a21oi_1
XFILLER_7_334 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1
+ net2302 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[136\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_98_639 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1 net3016 i_snitch.i_snitch_regfile.mem\[400\]
+ i_snitch.i_snitch_regfile.mem\[432\] i_snitch.i_snitch_regfile.mem\[464\] i_snitch.i_snitch_regfile.mem\[496\]
+ net2987 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0 net3001 i_snitch.i_snitch_regfile.mem\[391\]
+ i_snitch.i_snitch_regfile.mem\[423\] i_snitch.i_snitch_regfile.mem\[455\] i_snitch.i_snitch_regfile.mem\[487\]
+ net2974 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_79_886 VPWR VGND sg13g2_decap_8
XFILLER_78_330 VPWR VGND sg13g2_decap_8
XFILLER_66_525 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2777 net2912 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_38_205 VPWR VGND sg13g2_decap_8
XFILLER_38_216 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net89 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
XFILLER_94_889 VPWR VGND sg13g2_decap_8
XFILLER_93_366 VPWR VGND sg13g2_fill_2
XFILLER_47_772 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[3\]_sg13g2_a22oi_1_A1 uio_out_sg13g2_inv_1_Y_A shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_mux2_1_A1_1_X
+ cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 shift_reg_q\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_35_956 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2702 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_50_904 VPWR VGND sg13g2_decap_4
Xdata_pdata\[22\]_sg13g2_a21oi_1_A2 VGND VPWR net3162 data_pdata\[22\] data_pdata\[22\]_sg13g2_a21oi_1_A2_Y
+ net3154 sg13g2_a21oi_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ net2535 i_req_arb.data_i\[39\] i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2784
+ net2654 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ net2560 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
Xhold802 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net834 sg13g2_dlygate4sd3_1
Xhold813 i_snitch.i_snitch_regfile.mem\[47\] VPWR VGND net845 sg13g2_dlygate4sd3_1
Xhold835 i_snitch.i_snitch_regfile.mem\[53\] VPWR VGND net867 sg13g2_dlygate4sd3_1
Xhold824 i_snitch.i_snitch_regfile.mem\[454\] VPWR VGND net856 sg13g2_dlygate4sd3_1
Xhold846 i_snitch.i_snitch_regfile.mem\[486\] VPWR VGND net878 sg13g2_dlygate4sd3_1
XFILLER_104_928 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ net2602 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.wake_up_q\[1\] clknet_leaf_38_clk sg13g2_dfrbpq_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 net2518 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ net2755 VPWR VGND sg13g2_a22oi_1
Xhold868 i_snitch.i_snitch_regfile.mem\[72\] VPWR VGND net900 sg13g2_dlygate4sd3_1
Xhold857 data_pdata\[9\] VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold879 i_snitch.i_snitch_regfile.mem\[110\] VPWR VGND net911 sg13g2_dlygate4sd3_1
XFILLER_84_300 VPWR VGND sg13g2_decap_4
XFILLER_85_878 VPWR VGND sg13g2_decap_8
XFILLER_83_19 VPWR VGND sg13g2_fill_2
XFILLER_72_506 VPWR VGND sg13g2_fill_1
XFILLER_84_399 VPWR VGND sg13g2_fill_2
XFILLER_53_764 VPWR VGND sg13g2_decap_8
XFILLER_53_797 VPWR VGND sg13g2_fill_1
XFILLER_41_948 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[156\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1 net3016 i_snitch.i_snitch_regfile.mem\[402\]
+ i_snitch.i_snitch_regfile.mem\[434\] i_snitch.i_snitch_regfile.mem\[466\] i_snitch.i_snitch_regfile.mem\[498\]
+ net2987 i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_21_650 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y VGND VPWR net2520 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D
+ net1392 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B VPWR
+ VGND sg13g2_nand2_1
XFILLER_106_210 VPWR VGND sg13g2_decap_8
XFILLER_106_287 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ net77 VGND sg13g2_inv_1
XFILLER_57_20 VPWR VGND sg13g2_fill_2
XFILLER_0_576 VPWR VGND sg13g2_decap_8
XFILLER_91_804 VPWR VGND sg13g2_decap_4
XFILLER_75_388 VPWR VGND sg13g2_fill_1
XFILLER_29_783 VPWR VGND sg13g2_decap_8
Xdata_pdata\[6\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B net3154 data_pdata\[6\]_sg13g2_mux2_1_A0_X
+ data_pdata\[6\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A_sg13g2_o21ai_1_Y
+ net2528 VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A
+ VGND i_snitch.inst_addr_o\[13\] i_snitch.inst_addr_o\[14\] sg13g2_o21ai_1
XFILLER_43_263 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B
+ VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1 net3008 i_snitch.i_snitch_regfile.mem\[287\]
+ i_snitch.i_snitch_regfile.mem\[319\] i_snitch.i_snitch_regfile.mem\[351\] i_snitch.i_snitch_regfile.mem\[383\]
+ net2982 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2748 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A
+ sg13g2_or2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_nor3_1_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nor3_1
Xstrb_reg_q\[2\]_sg13g2_nor2_1_A net517 net2727 strb_reg_q\[2\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_99_937 VPWR VGND sg13g2_decap_8
XFILLER_98_436 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[426\]_sg13g2_a21o_1_A1 net3013 i_snitch.i_snitch_regfile.mem\[426\]
+ net2979 i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_a21o_1_A1_X VPWR VGND sg13g2_a21o_1
XFILLER_79_650 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ net2574 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[18\]_sg13g2_nor2_1_A net508 net2734 shift_reg_q\[18\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0 net3134 i_snitch.i_snitch_regfile.mem\[279\]
+ i_snitch.i_snitch_regfile.mem\[311\] i_snitch.i_snitch_regfile.mem\[343\] i_snitch.i_snitch_regfile.mem\[375\]
+ net3113 i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_66_377 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[176\] clknet_leaf_89_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[350\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C
+ VPWR VGND sg13g2_nor2_1
XFILLER_34_252 VPWR VGND sg13g2_fill_1
XFILLER_35_775 VPWR VGND sg13g2_fill_2
XFILLER_62_572 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y i_snitch.pc_d\[12\] i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2 net2308 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_50_767 VPWR VGND sg13g2_fill_1
XFILLER_23_959 VPWR VGND sg13g2_decap_4
XFILLER_33_1014 VPWR VGND sg13g2_decap_8
Xhold610 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\] VPWR
+ VGND net642 sg13g2_dlygate4sd3_1
Xhold621 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\] VPWR
+ VGND net653 sg13g2_dlygate4sd3_1
Xhold632 i_snitch.i_snitch_regfile.mem\[328\] VPWR VGND net664 sg13g2_dlygate4sd3_1
Xhold643 i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y VPWR VGND net675 sg13g2_dlygate4sd3_1
Xhold654 data_pdata\[2\] VPWR VGND net686 sg13g2_dlygate4sd3_1
XFILLER_103_224 VPWR VGND sg13g2_decap_8
Xhold676 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\] VPWR
+ VGND net708 sg13g2_dlygate4sd3_1
Xhold665 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\] VPWR
+ VGND net697 sg13g2_dlygate4sd3_1
Xhold687 data_pdata\[6\] VPWR VGND net719 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xhold698 data_pdata\[17\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net730 sg13g2_dlygate4sd3_1
XFILLER_100_931 VPWR VGND sg13g2_decap_8
XFILLER_97_491 VPWR VGND sg13g2_fill_1
Xhold1343 i_snitch.inst_addr_o\[13\] VPWR VGND net1375 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2375 net862 net2665 net2743 VPWR VGND sg13g2_a22oi_1
Xhold1332 i_snitch.i_snitch_regfile.mem\[99\] VPWR VGND net1364 sg13g2_dlygate4sd3_1
Xhold1321 i_snitch.i_snitch_regfile.mem\[101\] VPWR VGND net1353 sg13g2_dlygate4sd3_1
Xhold1310 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\] VPWR
+ VGND net1342 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0 net3130 i_snitch.i_snitch_regfile.mem\[398\]
+ i_snitch.i_snitch_regfile.mem\[430\] i_snitch.i_snitch_regfile.mem\[462\] i_snitch.i_snitch_regfile.mem\[494\]
+ net3109 i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold1354 i_snitch.inst_addr_o\[29\] VPWR VGND net1386 sg13g2_dlygate4sd3_1
Xhold1365 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[1\] VPWR VGND net1397 sg13g2_dlygate4sd3_1
Xhold1376 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q VPWR VGND net1408 sg13g2_dlygate4sd3_1
XFILLER_58_889 VPWR VGND sg13g2_fill_1
XFILLER_58_878 VPWR VGND sg13g2_decap_4
XFILLER_17_219 VPWR VGND sg13g2_fill_1
XFILLER_85_697 VPWR VGND sg13g2_fill_1
XFILLER_72_358 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q
+ net3229 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_53_561 VPWR VGND sg13g2_fill_2
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C net3163 i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nand2b_1_B_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y VGND VPWR data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D
+ sg13g2_nor4_2
XFILLER_80_380 VPWR VGND sg13g2_decap_8
XFILLER_43_55 VPWR VGND sg13g2_fill_2
Xdata_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2 data_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ net3070 net2714 data_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_40_244 VPWR VGND sg13g2_decap_4
XFILLER_41_756 VPWR VGND sg13g2_fill_2
XFILLER_22_970 VPWR VGND sg13g2_fill_2
XFILLER_40_299 VPWR VGND sg13g2_fill_2
Xdata_pdata\[26\]_sg13g2_mux2_1_A1 rsp_data_q\[26\] net818 net3048 data_pdata\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_104_0 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\] net2617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[196\] clknet_leaf_13_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[363\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[363\] net2807 sg13g2_o21ai_1
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_96_929 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A
+ net3087 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_B1
+ VPWR VGND net120 sg13g2_nand4_1
XFILLER_68_30 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[502\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_49_801 VPWR VGND sg13g2_decap_8
XFILLER_76_620 VPWR VGND sg13g2_decap_8
XFILLER_0_351 VPWR VGND sg13g2_decap_8
XFILLER_1_874 VPWR VGND sg13g2_decap_8
XFILLER_91_601 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_nor3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_76_675 VPWR VGND sg13g2_fill_1
XFILLER_76_664 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q net3310 VGND VPWR i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[44\] clknet_leaf_69_clk sg13g2_dfrbpq_1
XFILLER_76_697 VPWR VGND sg13g2_fill_1
XFILLER_56_1025 VPWR VGND sg13g2_decap_4
XFILLER_32_712 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2757 net2303
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2517 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_16_285 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_277 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A_Y i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_12_480 VPWR VGND sg13g2_decap_8
XFILLER_76_4 VPWR VGND sg13g2_fill_1
XFILLER_9_985 VPWR VGND sg13g2_decap_8
XFILLER_99_712 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[492\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[492\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net1112 net2691 net2857 VPWR VGND sg13g2_a22oi_1
XFILLER_98_211 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B
+ net93 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_98_244 VPWR VGND sg13g2_fill_2
XFILLER_59_609 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[19\]_sg13g2_a22oi_1_A1 shift_reg_q\[19\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ net3055 net3046 shift_reg_q\[19\] VPWR VGND sg13g2_a22oi_1
XFILLER_100_205 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1
+ VGND net96 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_86_417 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q
+ net3229 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
XFILLER_104_28 VPWR VGND sg13g2_decap_8
XFILLER_95_973 VPWR VGND sg13g2_decap_8
XFILLER_55_815 VPWR VGND sg13g2_fill_1
XFILLER_81_100 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A_Y net3031 sg13g2_o21ai_1
XFILLER_39_388 VPWR VGND sg13g2_decap_8
XFILLER_82_678 VPWR VGND sg13g2_decap_4
XFILLER_82_667 VPWR VGND sg13g2_fill_2
XFILLER_70_829 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2560 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_82_689 VPWR VGND sg13g2_decap_4
XFILLER_81_177 VPWR VGND sg13g2_decap_4
XFILLER_81_166 VPWR VGND sg13g2_fill_1
XFILLER_35_572 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2572 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ net2538 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2758 net2304
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1 net2518 sg13g2_a221oi_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y net414 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C
+ net2519 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1 VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1
+ net95 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ net2719 i_req_arb.data_i\[38\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[311\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[311\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2647 net2780 net2318 net1182 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_C i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_B1
+ i_snitch.inst_addr_o\[17\] net2313 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2 VPWR
+ VGND sg13g2_and3_1
Xfanout3309 net3311 net3309 VPWR VGND sg13g2_buf_8
Xfanout2608 net2608 net2609 VPWR VGND sg13g2_buf_16
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q net3257 VGND VPWR i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[64\] clknet_leaf_49_clk sg13g2_dfrbpq_1
Xhold440 strb_reg_q\[4\] VPWR VGND net472 sg13g2_dlygate4sd3_1
XFILLER_8_7 VPWR VGND sg13g2_decap_8
Xhold451 shift_reg_q\[21\] VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold462 i_snitch.i_snitch_regfile.mem\[97\] VPWR VGND net494 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2358
+ sg13g2_o21ai_1
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_2_649 VPWR VGND sg13g2_decap_8
Xhold484 shift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net516 sg13g2_dlygate4sd3_1
Xhold473 i_snitch.i_snitch_regfile.mem\[257\] VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold495 shift_reg_q\[0\] VPWR VGND net527 sg13g2_dlygate4sd3_1
Xfanout2619 net2620 net2619 VPWR VGND sg13g2_buf_8
XFILLER_86_951 VPWR VGND sg13g2_decap_8
Xhold1151 rsp_data_q\[8\] VPWR VGND net1183 sg13g2_dlygate4sd3_1
XFILLER_79_1014 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[312\]
+ net3022 i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_a21oi_1_A1_Y net2990 sg13g2_a21oi_1
Xhold1140 i_snitch.i_snitch_regfile.mem\[121\] VPWR VGND net1172 sg13g2_dlygate4sd3_1
XFILLER_46_848 VPWR VGND sg13g2_fill_1
Xhold1173 i_snitch.i_snitch_regfile.mem\[314\] VPWR VGND net1205 sg13g2_dlygate4sd3_1
Xhold1184 i_snitch.i_snitch_regfile.mem\[126\] VPWR VGND net1216 sg13g2_dlygate4sd3_1
Xhold1162 i_snitch.i_snitch_regfile.mem\[366\] VPWR VGND net1194 sg13g2_dlygate4sd3_1
Xhold1195 rsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1227
+ sg13g2_dlygate4sd3_1
XFILLER_33_509 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3062 net1347 net3063 rsp_data_q\[21\] VPWR VGND sg13g2_a22oi_1
XFILLER_54_870 VPWR VGND sg13g2_fill_1
XFILLER_54_54 VPWR VGND sg13g2_decap_4
XFILLER_26_561 VPWR VGND sg13g2_fill_2
XFILLER_60_339 VPWR VGND sg13g2_decap_8
XFILLER_9_215 VPWR VGND sg13g2_decap_8
XFILLER_16_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_103_1012 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2429 i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_A1 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_86_1007 VPWR VGND sg13g2_decap_8
Xclkload29 clknet_leaf_31_clk clkload29/X VPWR VGND sg13g2_buf_8
Xclkload18 clkload18/Y clknet_leaf_27_clk VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_dfrbpq_1_Q_D VGND net2400 net310
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B
+ VGND net2745 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
XFILLER_6_977 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_68_428 VPWR VGND sg13g2_fill_2
XFILLER_1_671 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xdata_pdata\[5\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net677 data_pdata\[5\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y_sg13g2_nor3_1_A i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[29\]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A_Y i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nor3_2
XFILLER_77_984 VPWR VGND sg13g2_decap_8
XFILLER_48_130 VPWR VGND sg13g2_fill_2
XFILLER_37_804 VPWR VGND sg13g2_fill_1
XFILLER_92_976 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp
+ net91 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X VPWR VGND
+ sg13g2_and2_1
XFILLER_52_829 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[331\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2404 net709 net2680 net2797 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_nand2_1_A_Y net3028 net2997 i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]
+ net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_2
Xi_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[84\] clknet_leaf_60_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nor2_1_B
+ net2565 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1
+ net873 net655 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.data_o\[39\]_sg13g2_o21ai_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2496 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_105_308 VPWR VGND sg13g2_decap_8
XFILLER_87_704 VPWR VGND sg13g2_fill_2
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C
+ net2924 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B
+ net2927 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C_Y
+ VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ sg13g2_nand4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_101_503 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor3_2
XFILLER_8_1018 VPWR VGND sg13g2_decap_8
XFILLER_87_748 VPWR VGND sg13g2_decap_4
XFILLER_83_921 VPWR VGND sg13g2_decap_8
XFILLER_27_325 VPWR VGND sg13g2_decap_4
XFILLER_82_442 VPWR VGND sg13g2_fill_1
Xstate_sg13g2_dfrbpq_1_Q net3184 VGND VPWR state_sg13g2_dfrbpq_1_Q_D state clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_83_998 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND net2557 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_24_68 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net89 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2366
+ sg13g2_o21ai_1
Xfanout3117 net3118 net3117 VPWR VGND sg13g2_buf_8
Xfanout3106 net3107 net3106 VPWR VGND sg13g2_buf_8
Xfanout3128 net3128 net3132 VPWR VGND sg13g2_buf_16
Xfanout3139 net3140 net3139 VPWR VGND sg13g2_buf_8
XFILLER_3_969 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2460 net2739 i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
Xfanout2405 net2406 net2405 VPWR VGND sg13g2_buf_8
Xfanout2416 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2416 VPWR VGND sg13g2_buf_1
XFILLER_105_875 VPWR VGND sg13g2_decap_8
Xfanout2427 net2428 net2427 VPWR VGND sg13g2_buf_8
Xfanout2449 net2450 net2449 VPWR VGND sg13g2_buf_8
Xfanout2438 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2438 VPWR
+ VGND sg13g2_buf_8
XFILLER_104_385 VPWR VGND sg13g2_decap_8
XFILLER_78_748 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N
+ sg13g2_a21oi_2
XFILLER_93_729 VPWR VGND sg13g2_decap_8
XFILLER_93_718 VPWR VGND sg13g2_fill_1
XFILLER_77_258 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[351\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2403 net813 net2645 net2796 VPWR VGND sg13g2_a22oi_1
XFILLER_1_28 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B net2817
+ i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_65_42 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_18_369 VPWR VGND sg13g2_decap_8
XFILLER_92_1011 VPWR VGND sg13g2_decap_8
XFILLER_61_648 VPWR VGND sg13g2_decap_4
XFILLER_60_136 VPWR VGND sg13g2_fill_1
XFILLER_26_380 VPWR VGND sg13g2_fill_2
XFILLER_42_840 VPWR VGND sg13g2_decap_8
XFILLER_53_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[352\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[352\]
+ net3124 i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_a21oi_1_A1_Y net2941 sg13g2_a21oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2590 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2584 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_mux4_1_X
+ net3123 i_snitch.sb_q\[8\] i_snitch.sb_q\[9\] i_snitch.sb_q\[10\] i_snitch.sb_q\[11\]
+ net3103 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux4_1
XFILLER_60_7 VPWR VGND sg13g2_fill_1
XFILLER_96_512 VPWR VGND sg13g2_decap_8
XFILLER_69_737 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net3039 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2
+ net2504 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_96_523 VPWR VGND sg13g2_fill_2
Xfanout2972 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2972 VPWR VGND sg13g2_buf_8
Xfanout2961 net2962 net2961 VPWR VGND sg13g2_buf_8
Xfanout2950 net2951 net2950 VPWR VGND sg13g2_buf_8
XFILLER_83_206 VPWR VGND sg13g2_fill_1
Xfanout2983 net2984 net2983 VPWR VGND sg13g2_buf_8
Xfanout2994 net2995 net2994 VPWR VGND sg13g2_buf_8
XFILLER_77_792 VPWR VGND sg13g2_fill_2
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_92_762 VPWR VGND sg13g2_decap_8
XFILLER_92_740 VPWR VGND sg13g2_fill_1
XFILLER_25_807 VPWR VGND sg13g2_decap_8
XFILLER_80_924 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q
+ net3198 VGND VPWR net585 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
XFILLER_33_884 VPWR VGND sg13g2_fill_1
XFILLER_20_567 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ net95 i_req_arb.data_i\[39\] i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ net2719 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[371\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net988 net2469 net2271 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1_A2
+ net2940 net3120 VPWR VGND sg13g2_nand2_1
XFILLER_105_105 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1
+ net2489 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C
+ VPWR VGND sg13g2_and3_1
Xtarget_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B_Y
+ VPWR VGND net3164 sg13g2_nand3b_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[0\] net747 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_99_372 VPWR VGND sg13g2_decap_8
XFILLER_102_856 VPWR VGND sg13g2_decap_8
XFILLER_101_322 VPWR VGND sg13g2_decap_8
XFILLER_87_567 VPWR VGND sg13g2_fill_1
XFILLER_74_239 VPWR VGND sg13g2_fill_1
XFILLER_68_770 VPWR VGND sg13g2_decap_4
XFILLER_83_751 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B
+ net2834 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ net2981 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[372\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[372\]
+ net3137 i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
XFILLER_55_453 VPWR VGND sg13g2_decap_8
XFILLER_16_807 VPWR VGND sg13g2_fill_2
XFILLER_82_250 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N_Y
+ net3176 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_55_464 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[506\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2254 net2367 net1136 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y
+ VPWR VGND sg13g2_inv_2
XFILLER_24_895 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[401\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_51_77 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1198 net2456 net2262 VPWR VGND sg13g2_a22oi_1
XFILLER_100_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[450\]_sg13g2_nor3_1_A net1270 net2739 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2722 i_snitch.inst_addr_o\[10\] sg13g2_a21oi_2
XFILLER_3_700 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A
+ net3074 net2537 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_mux2_1_A1
+ net854 net561 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_2_232 VPWR VGND sg13g2_fill_1
XFILLER_105_694 VPWR VGND sg13g2_fill_1
XFILLER_104_182 VPWR VGND sg13g2_decap_8
XFILLER_78_534 VPWR VGND sg13g2_decap_4
Xfanout2257 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2257 VPWR VGND sg13g2_buf_8
Xfanout2246 net2247 net2246 VPWR VGND sg13g2_buf_8
Xfanout2268 net2269 net2268 VPWR VGND sg13g2_buf_8
Xfanout2279 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y
+ net2279 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR net429 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_93_537 VPWR VGND sg13g2_decap_8
XFILLER_19_645 VPWR VGND sg13g2_fill_2
XFILLER_19_667 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_q\[7\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.sb_d\[7\] i_snitch.sb_q\[7\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_61_401 VPWR VGND sg13g2_decap_4
XFILLER_73_294 VPWR VGND sg13g2_decap_4
XFILLER_62_968 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2285 net2387 net1317 VPWR VGND sg13g2_a22oi_1
XFILLER_21_309 VPWR VGND sg13g2_fill_2
XFILLER_61_489 VPWR VGND sg13g2_fill_1
XFILLER_14_372 VPWR VGND sg13g2_decap_4
XFILLER_30_832 VPWR VGND sg13g2_decap_4
XFILLER_42_692 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2779
+ net2656 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ net2429 VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2489 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ sg13g2_o21ai_1
XFILLER_102_119 VPWR VGND sg13g2_decap_8
XFILLER_97_887 VPWR VGND sg13g2_decap_8
XFILLER_57_707 VPWR VGND sg13g2_fill_2
Xfanout2780 net2781 net2780 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[82\] net2987 VPWR VGND sg13g2_nand2_1
XFILLER_99_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_60 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2794 net2906 i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_38_932 VPWR VGND sg13g2_fill_1
Xfanout2791 net2792 net2791 VPWR VGND sg13g2_buf_8
XFILLER_49_280 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2733 shift_reg_q\[22\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[18\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[18\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[419\]_sg13g2_nor3_1_A net1301 net2860 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[421\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[210\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net968 net2441 net2272 VPWR VGND sg13g2_a22oi_1
XFILLER_53_979 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2530 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_191 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2872
+ net2673 VPWR VGND sg13g2_nand2_1
XFILLER_82_1021 VPWR VGND sg13g2_decap_8
XFILLER_88_854 VPWR VGND sg13g2_decap_8
XFILLER_0_758 VPWR VGND sg13g2_decap_8
XFILLER_87_386 VPWR VGND sg13g2_decap_4
XFILLER_75_537 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[101\]
+ net2800 sg13g2_o21ai_1
XFILLER_101_196 VPWR VGND sg13g2_decap_8
XFILLER_75_559 VPWR VGND sg13g2_fill_2
XFILLER_56_740 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1
+ net2748 net2579 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[341\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2658 VPWR VGND sg13g2_nand2_1
XFILLER_16_604 VPWR VGND sg13g2_fill_2
XFILLER_28_475 VPWR VGND sg13g2_decap_8
XFILLER_29_987 VPWR VGND sg13g2_fill_1
XFILLER_71_743 VPWR VGND sg13g2_fill_1
XFILLER_71_732 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B
+ net115 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a21o_1
XFILLER_15_158 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3040
+ net2667 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[104\]
+ net2998 i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2774
+ net2693 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[88\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net766 net2666 net2787 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A_Y net2846 i_snitch.i_snitch_regfile.mem\[343\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[441\] clknet_leaf_114_clk sg13g2_dfrbpq_1
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_79_854 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[230\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net918 net2900 net2876 VPWR VGND sg13g2_a22oi_1
XFILLER_94_868 VPWR VGND sg13g2_decap_8
XFILLER_19_420 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X
+ VPWR VGND sg13g2_and4_1
XFILLER_59_1001 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B_sg13g2_inv_1_Y
+ VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2676 VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1271 net3063 rsp_data_q\[19\] VPWR VGND sg13g2_a22oi_1
XFILLER_62_765 VPWR VGND sg13g2_fill_1
XFILLER_61_253 VPWR VGND sg13g2_fill_2
XFILLER_50_927 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[89\]
+ net2840 i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
XFILLER_22_618 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A
+ sg13g2_or2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR net707 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
Xdata_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[9\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[25\]_sg13g2_nand2b_1_B_Y net3149 data_pdata\[17\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[9\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
Xhold803 i_snitch.i_snitch_regfile.mem\[238\] VPWR VGND net835 sg13g2_dlygate4sd3_1
Xhold836 i_snitch.i_snitch_regfile.mem\[504\] VPWR VGND net868 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2878
+ net2660 VPWR VGND sg13g2_nand2_1
Xhold825 i_snitch.i_snitch_regfile.mem\[217\] VPWR VGND net857 sg13g2_dlygate4sd3_1
Xhold814 data_pdata\[29\] VPWR VGND net846 sg13g2_dlygate4sd3_1
XFILLER_104_907 VPWR VGND sg13g2_decap_8
XFILLER_103_406 VPWR VGND sg13g2_decap_8
XFILLER_89_618 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q_sg13g2_dfrbpq_1_Q net3252 VGND VPWR
+ i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2991 net2852 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2
+ net2629 sg13g2_a21oi_1
XFILLER_66_1027 VPWR VGND sg13g2_fill_2
Xhold847 i_snitch.i_snitch_regfile.mem\[344\] VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold869 data_pdata\[12\] VPWR VGND net901 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B
+ net2639 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
Xhold858 data_pdata\[9\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net890 sg13g2_dlygate4sd3_1
XFILLER_103_428 VPWR VGND sg13g2_fill_1
XFILLER_69_320 VPWR VGND sg13g2_fill_2
XFILLER_97_651 VPWR VGND sg13g2_fill_2
XFILLER_97_673 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[22\]_sg13g2_dfrbpq_1_Q net3231 VGND VPWR rsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[22\] clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_85_857 VPWR VGND sg13g2_decap_8
XFILLER_84_323 VPWR VGND sg13g2_decap_8
XFILLER_29_239 VPWR VGND sg13g2_decap_8
XFILLER_84_356 VPWR VGND sg13g2_decap_8
XFILLER_38_773 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_A1
+ net1386 VGND sg13g2_inv_1
XFILLER_80_551 VPWR VGND sg13g2_decap_8
XFILLER_80_540 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0 net3129 i_snitch.i_snitch_regfile.mem\[400\]
+ i_snitch.i_snitch_regfile.mem\[432\] i_snitch.i_snitch_regfile.mem\[464\] i_snitch.i_snitch_regfile.mem\[496\]
+ net3108 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_80_573 VPWR VGND sg13g2_decap_8
XFILLER_13_618 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[117\]
+ net2948 i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[461\] clknet_leaf_88_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[250\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net993 net2436 net2254 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nor3_1_A net1333 net2783 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
XFILLER_106_266 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2440
+ net2513 net2901 net2791 VPWR VGND sg13g2_a22oi_1
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_103_984 VPWR VGND sg13g2_decap_8
XFILLER_76_813 VPWR VGND sg13g2_fill_1
XFILLER_57_98 VPWR VGND sg13g2_decap_4
XFILLER_91_849 VPWR VGND sg13g2_decap_8
XFILLER_56_592 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR net613 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_43_242 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[444\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_8_600 VPWR VGND sg13g2_decap_4
XFILLER_11_150 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2462 VPWR VGND sg13g2_nand2_1
XFILLER_8_666 VPWR VGND sg13g2_decap_4
Xi_req_register.data_o\[38\]_sg13g2_mux2_1_X i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[38\] net3164 i_req_register.data_o\[38\]
+ VPWR VGND sg13g2_mux2_1
XFILLER_99_916 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2596 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[187\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_409 VPWR VGND sg13g2_fill_1
XFILLER_94_610 VPWR VGND sg13g2_fill_1
XFILLER_79_695 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_1 net3101 VPWR i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[97\] net2951 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[109\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_39_504 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2766
+ net2656 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[481\] clknet_leaf_75_clk sg13g2_dfrbpq_1
Xdata_pdata\[24\]_sg13g2_nand2b_1_B data_pdata\[24\]_sg13g2_nand2b_1_B_Y data_pdata\[24\]
+ net3159 VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_882 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net940 net2687 net2895 VPWR VGND sg13g2_a22oi_1
XFILLER_97_0 VPWR VGND sg13g2_decap_8
Xhold611 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\] VPWR
+ VGND net643 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xhold600 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\] VPWR
+ VGND net632 sg13g2_dlygate4sd3_1
XFILLER_104_704 VPWR VGND sg13g2_fill_1
Xhold633 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\] VPWR
+ VGND net665 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2551 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
Xhold622 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net654 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[271\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[271\]
+ net3029 i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_a21oi_1_A1_Y net2990 sg13g2_a21oi_1
Xhold644 data_pdata\[5\] VPWR VGND net676 sg13g2_dlygate4sd3_1
XFILLER_104_748 VPWR VGND sg13g2_fill_1
XFILLER_103_203 VPWR VGND sg13g2_decap_8
Xhold666 data_pdata\[4\] VPWR VGND net698 sg13g2_dlygate4sd3_1
Xhold677 i_snitch.i_snitch_regfile.mem\[331\] VPWR VGND net709 sg13g2_dlygate4sd3_1
Xhold688 data_pdata\[6\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net720 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[6\]
+ VGND net2293 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold655 data_pdata\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net687 sg13g2_dlygate4sd3_1
XFILLER_89_459 VPWR VGND sg13g2_fill_1
Xhold699 i_snitch.i_snitch_regfile.mem\[95\] VPWR VGND net731 sg13g2_dlygate4sd3_1
Xdata_pdata\[23\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net722 data_pdata\[23\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2466 net2268 net2387 net1220 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2592 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_100_910 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y net2309 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2 VPWR VGND sg13g2_nor2_1
XFILLER_76_109 VPWR VGND sg13g2_fill_1
Xhold1300 i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp
+ VPWR VGND net1332 sg13g2_dlygate4sd3_1
Xhold1333 rsp_data_q\[5\] VPWR VGND net1365 sg13g2_dlygate4sd3_1
XFILLER_85_632 VPWR VGND sg13g2_fill_2
Xhold1311 rsp_data_q\[9\] VPWR VGND net1343 sg13g2_dlygate4sd3_1
Xhold1322 rsp_data_q\[0\] VPWR VGND net1354 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2458 VPWR VGND sg13g2_nand2_1
XFILLER_40_1019 VPWR VGND sg13g2_decap_8
XFILLER_100_987 VPWR VGND sg13g2_decap_8
Xhold1377 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]
+ VPWR VGND net1409 sg13g2_dlygate4sd3_1
Xhold1366 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_A VPWR VGND net1398 sg13g2_dlygate4sd3_1
Xhold1344 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] VPWR
+ VGND net1376 sg13g2_dlygate4sd3_1
Xhold1355 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\] VPWR
+ VGND net1387 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[300\] clknet_leaf_69_clk sg13g2_dfrbpq_1
XFILLER_66_890 VPWR VGND sg13g2_fill_2
XFILLER_14_905 VPWR VGND sg13g2_decap_8
XFILLER_27_79 VPWR VGND sg13g2_fill_1
XFILLER_81_893 VPWR VGND sg13g2_decap_8
XFILLER_41_713 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[406\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[406\]
+ net3030 i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_a21oi_1_A1_Y net2992 sg13g2_a21oi_1
XFILLER_53_595 VPWR VGND sg13g2_decap_8
XFILLER_43_45 VPWR VGND sg13g2_fill_1
XFILLER_40_223 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ VGND i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[129\] clknet_leaf_75_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2783
+ net2658 VPWR VGND sg13g2_nand2_1
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_96_908 VPWR VGND sg13g2_decap_8
XFILLER_1_853 VPWR VGND sg13g2_decap_8
XFILLER_89_993 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_a21o_1_A1 net3123 i_snitch.i_snitch_regfile.mem\[511\]
+ net2941 i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_a21o_1_A1_X VPWR VGND sg13g2_a21o_1
XFILLER_103_781 VPWR VGND sg13g2_decap_8
XFILLER_102_280 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2551 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y
+ VGND VPWR net2704 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VGND net2589 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_64_827 VPWR VGND sg13g2_decap_4
XFILLER_91_679 VPWR VGND sg13g2_fill_1
XFILLER_44_562 VPWR VGND sg13g2_decap_8
XFILLER_32_702 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_7 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net451 net2405 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net2429 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2
+ net2493 net533 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0 net3024 i_snitch.i_snitch_regfile.mem\[407\]
+ i_snitch.i_snitch_regfile.mem\[439\] i_snitch.i_snitch_regfile.mem\[471\] i_snitch.i_snitch_regfile.mem\[503\]
+ net2991 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_13_960 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2627 net2851 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2328
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[425\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2384 net779 net2685 net2861 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q net3255 VGND VPWR i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[320\] clknet_leaf_17_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2700 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_86_429 VPWR VGND sg13g2_decap_8
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_95_952 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2b_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_nor2_1_B
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_67_621 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[417\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net524 net2381 VPWR VGND sg13g2_nand2_1
XFILLER_39_334 VPWR VGND sg13g2_fill_1
XFILLER_82_602 VPWR VGND sg13g2_fill_1
Xdata_pdata\[30\]_sg13g2_mux2_1_A1 rsp_data_q\[30\] net1054 net3050 data_pdata\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_66_186 VPWR VGND sg13g2_fill_2
XFILLER_23_724 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y
+ net2750 VPWR VGND net86 sg13g2_nand2b_2
Xrsp_data_ready_sg13g2_nor2b_1_Y net914 net2 rsp_data_ready VPWR VGND sg13g2_nor2b_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[149\] clknet_leaf_98_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[455\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[455\] net2947 VPWR VGND sg13g2_nand2_1
XFILLER_23_735 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y net2954
+ i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xfanout2609 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N_Y
+ net2609 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2759 net2304
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2517 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
Xhold430 shift_reg_q\[15\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net462 sg13g2_dlygate4sd3_1
Xhold441 strb_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net473 sg13g2_dlygate4sd3_1
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_2_628 VPWR VGND sg13g2_decap_8
Xhold452 shift_reg_q\[21\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold463 i_snitch.i_snitch_regfile.mem\[385\] VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold474 shift_reg_q\[6\] VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold485 strb_reg_q\[2\] VPWR VGND net517 sg13g2_dlygate4sd3_1
Xhold496 shift_reg_q\[0\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net528 sg13g2_dlygate4sd3_1
XFILLER_104_578 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[346\] VGND sg13g2_inv_1
XFILLER_86_930 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2348
+ sg13g2_o21ai_1
XFILLER_58_621 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_740 VPWR VGND sg13g2_decap_8
XFILLER_85_462 VPWR VGND sg13g2_fill_1
Xhold1141 i_snitch.i_snitch_regfile.mem\[380\] VPWR VGND net1173 sg13g2_dlygate4sd3_1
Xhold1130 i_snitch.i_snitch_regfile.mem\[315\] VPWR VGND net1162 sg13g2_dlygate4sd3_1
XFILLER_100_784 VPWR VGND sg13g2_decap_8
Xhold1152 rsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1184 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X
+ VPWR VGND sg13g2_or3_1
Xhold1163 i_snitch.i_snitch_regfile.mem\[308\] VPWR VGND net1195 sg13g2_dlygate4sd3_1
XFILLER_57_164 VPWR VGND sg13g2_decap_8
Xhold1185 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\] VPWR
+ VGND net1217 sg13g2_dlygate4sd3_1
Xshift_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2733 shift_reg_q\[10\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[6\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_45_315 VPWR VGND sg13g2_fill_1
Xhold1174 i_snitch.i_snitch_regfile.mem\[355\] VPWR VGND net1206 sg13g2_dlygate4sd3_1
Xhold1196 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\] VPWR
+ VGND net1228 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2464 net2250 net2381 net1214 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2
+ net3179 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_14_779 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q net3315 VGND VPWR i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[340\] clknet_leaf_66_clk sg13g2_dfrbpq_1
XFILLER_13_289 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1_sg13g2_mux2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]
+ net3182 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2392
+ sg13g2_o21ai_1
Xclkload19 VPWR clkload19/Y clknet_leaf_30_clk VGND sg13g2_inv_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1
+ VPWR VGND i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A_Y
+ i_snitch.inst_addr_o\[24\] i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N_B
+ net2525 sg13g2_a221oi_1
XFILLER_6_956 VPWR VGND sg13g2_decap_8
XFILLER_96_705 VPWR VGND sg13g2_fill_2
XFILLER_95_215 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2
+ VPWR VGND sg13g2_and4_1
XFILLER_1_650 VPWR VGND sg13g2_decap_8
XFILLER_89_790 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y
+ i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[169\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_23_1025 VPWR VGND sg13g2_decap_4
XFILLER_91_410 VPWR VGND sg13g2_decap_8
XFILLER_92_955 VPWR VGND sg13g2_decap_8
XFILLER_63_145 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2833
+ VPWR i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_1_Y
+ sg13g2_o21ai_1
XFILLER_48_197 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2478 i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2471 net2879 i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
XFILLER_91_476 VPWR VGND sg13g2_fill_1
XFILLER_45_882 VPWR VGND sg13g2_fill_1
XFILLER_17_551 VPWR VGND sg13g2_fill_2
XFILLER_60_885 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ net2684 net2747 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A net45
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2937 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ net2932 sg13g2_a21oi_1
XFILLER_9_772 VPWR VGND sg13g2_decap_8
XFILLER_9_761 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0_X
+ net2938 net2931 i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_99_532 VPWR VGND sg13g2_fill_2
XFILLER_5_60 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[476\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y
+ VGND VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B
+ sg13g2_nor4_2
XFILLER_59_418 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[465\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[465\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net774 net2663 net2741 VPWR VGND sg13g2_a22oi_1
XFILLER_83_900 VPWR VGND sg13g2_decap_8
XFILLER_95_793 VPWR VGND sg13g2_decap_8
XFILLER_95_771 VPWR VGND sg13g2_fill_1
XFILLER_83_977 VPWR VGND sg13g2_decap_8
XFILLER_82_432 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[360\] clknet_leaf_74_clk sg13g2_dfrbpq_1
XFILLER_82_465 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2419 sg13g2_a21oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A
+ net123 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xrsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1384 net3063 net1349 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2334
+ sg13g2_o21ai_1
XFILLER_10_204 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[189\] clknet_leaf_96_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ net2549 VGND sg13g2_inv_1
Xfanout3129 net3131 net3129 VPWR VGND sg13g2_buf_8
Xfanout3118 net3121 net3118 VPWR VGND sg13g2_buf_8
Xfanout3107 net3110 net3107 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[356\]_sg13g2_o21ai_1_A1 net2969 VPWR i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[356\] net2803 sg13g2_o21ai_1
XFILLER_105_854 VPWR VGND sg13g2_decap_8
Xfanout2417 net2418 net2417 VPWR VGND sg13g2_buf_2
XFILLER_3_948 VPWR VGND sg13g2_decap_8
Xfanout2406 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2406 VPWR VGND sg13g2_buf_8
XFILLER_104_364 VPWR VGND sg13g2_decap_8
Xfanout2428 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A_X
+ net2428 VPWR VGND sg13g2_buf_8
Xfanout2439 net2441 net2439 VPWR VGND sg13g2_buf_8
XFILLER_93_708 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[37\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[37\] clknet_leaf_108_clk sg13g2_dfrbpq_1
Xi_snitch.inst_addr_o\[20\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.pc_d\[20\]
+ i_snitch.inst_addr_o\[20\] clknet_leaf_52_clk sg13g2_dfrbpq_2
XFILLER_18_304 VPWR VGND sg13g2_fill_2
XFILLER_74_955 VPWR VGND sg13g2_decap_4
XFILLER_73_498 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_119_clk clknet_5_1__leaf_clk clknet_leaf_119_clk VPWR VGND sg13g2_buf_8
XFILLER_60_159 VPWR VGND sg13g2_fill_2
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_5_296 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[380\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_69_749 VPWR VGND sg13g2_decap_8
Xfanout2962 net2967 net2962 VPWR VGND sg13g2_buf_8
Xfanout2940 net2941 net2940 VPWR VGND sg13g2_buf_8
Xfanout2973 net2976 net2973 VPWR VGND sg13g2_buf_8
XFILLER_2_992 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q
+ net3191 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
Xfanout2951 net2953 net2951 VPWR VGND sg13g2_buf_8
XFILLER_77_760 VPWR VGND sg13g2_fill_2
Xfanout2984 net2996 net2984 VPWR VGND sg13g2_buf_8
Xfanout2995 net2996 net2995 VPWR VGND sg13g2_buf_8
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
XFILLER_76_292 VPWR VGND sg13g2_fill_2
XFILLER_65_955 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y net710 VPWR i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1
+ VGND i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D
+ sg13g2_o21ai_1
XFILLER_92_796 VPWR VGND sg13g2_fill_2
XFILLER_80_903 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A_Y net2982 i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net3027 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2363
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_B_sg13g2_nand2_1_Y i_snitch.pc_d\[22\]_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_B2 net2308 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[332\] VGND sg13g2_inv_1
XFILLER_51_104 VPWR VGND sg13g2_fill_2
XFILLER_17_370 VPWR VGND sg13g2_decap_8
XFILLER_33_830 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[376\]_sg13g2_o21ai_1_A1 net2972 VPWR i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[376\] net2806 sg13g2_o21ai_1
XFILLER_33_852 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_32_395 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2431 net2263 net2317 net1243 VPWR VGND sg13g2_a22oi_1
XFILLER_106_607 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1 VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_106_618 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q net3215 VGND VPWR i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[57\] clknet_leaf_113_clk sg13g2_dfrbpq_1
XFILLER_99_351 VPWR VGND sg13g2_decap_8
XFILLER_87_502 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2511 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_102_835 VPWR VGND sg13g2_decap_8
XFILLER_101_301 VPWR VGND sg13g2_decap_8
XFILLER_99_395 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.inst_addr_o\[24\]
+ net2525 VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[305\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[305\]
+ net3020 i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_a21oi_1_A1_Y net2992 sg13g2_a21oi_1
XFILLER_19_36 VPWR VGND sg13g2_fill_1
XFILLER_101_389 VPWR VGND sg13g2_fill_1
XFILLER_101_378 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_A1
+ net2306 i_snitch.pc_d\[19\] i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
XFILLER_76_1018 VPWR VGND sg13g2_decap_8
XFILLER_82_284 VPWR VGND sg13g2_fill_1
XFILLER_43_627 VPWR VGND sg13g2_decap_4
XFILLER_11_524 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
XFILLER_23_395 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y net558 VPWR i_snitch.sb_d\[13\] VGND net2292
+ i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_7_539 VPWR VGND sg13g2_decap_8
XFILLER_13_1013 VPWR VGND sg13g2_decap_8
XFILLER_104_161 VPWR VGND sg13g2_decap_8
Xfanout2258 net2259 net2258 VPWR VGND sg13g2_buf_8
Xfanout2247 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ net2247 VPWR VGND sg13g2_buf_8
Xfanout2269 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ net2269 VPWR VGND sg13g2_buf_8
XFILLER_93_516 VPWR VGND sg13g2_decap_8
XFILLER_65_229 VPWR VGND sg13g2_fill_1
XFILLER_65_207 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2418 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_18_112 VPWR VGND sg13g2_fill_1
XFILLER_46_454 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[462\] VGND sg13g2_inv_1
XFILLER_15_863 VPWR VGND sg13g2_fill_2
XFILLER_70_980 VPWR VGND sg13g2_fill_2
XFILLER_14_351 VPWR VGND sg13g2_fill_1
XFILLER_25_90 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[77\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_42_671 VPWR VGND sg13g2_decap_8
XFILLER_41_170 VPWR VGND sg13g2_decap_4
XFILLER_30_888 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ net2583 VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VGND net2594 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D
+ sg13g2_nand4_1
XFILLER_6_572 VPWR VGND sg13g2_fill_1
Xdata_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2 data_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ net3070 net2714 data_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2593 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ net2587 sg13g2_a21oi_1
XFILLER_96_321 VPWR VGND sg13g2_decap_8
XFILLER_97_866 VPWR VGND sg13g2_decap_8
XFILLER_96_354 VPWR VGND sg13g2_fill_2
XFILLER_96_332 VPWR VGND sg13g2_fill_2
Xfanout2781 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X
+ net2781 VPWR VGND sg13g2_buf_8
Xfanout2770 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2_X
+ net2770 VPWR VGND sg13g2_buf_8
XFILLER_99_1007 VPWR VGND sg13g2_decap_8
Xfanout2792 net2793 net2792 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_Y
+ net2744 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ net95 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X
+ VPWR VGND sg13g2_or4_1
XFILLER_77_590 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y VPWR
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ net2626 sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_52_402 VPWR VGND sg13g2_fill_1
Xdata_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C i_snitch.i_snitch_lsu.metadata_q\[1\]
+ data_pdata\[19\]_sg13g2_mux2_1_A0_X data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y
+ VPWR VGND net3150 sg13g2_nand3b_1
XFILLER_92_571 VPWR VGND sg13g2_fill_1
XFILLER_53_936 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y net3135 sg13g2_o21ai_1
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_25_638 VPWR VGND sg13g2_fill_2
XFILLER_21_822 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net2429 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2
+ net2493 net820 VPWR VGND sg13g2_a22oi_1
XFILLER_106_448 VPWR VGND sg13g2_fill_2
XFILLER_82_1000 VPWR VGND sg13g2_decap_8
XFILLER_87_321 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_a22oi_1_B2_Y
+ net2404 net879 net2666 net2797 VPWR VGND sg13g2_a22oi_1
XFILLER_0_737 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.gpr_waddr\[5\] data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nand2_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_75_516 VPWR VGND sg13g2_decap_8
XFILLER_101_175 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C net2312 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.inst_addr_o\[1\] i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_B1 VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[97\] clknet_leaf_104_clk sg13g2_dfrbpq_1
XFILLER_28_421 VPWR VGND sg13g2_decap_4
XFILLER_29_933 VPWR VGND sg13g2_decap_8
XFILLER_56_785 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ VGND i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_56_796 VPWR VGND sg13g2_fill_1
XFILLER_70_243 VPWR VGND sg13g2_fill_2
XFILLER_102_84 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_50_clk clknet_5_24__leaf_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_8_815 VPWR VGND sg13g2_fill_2
XFILLER_12_877 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[3\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR rsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[3\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_7_39 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2870
+ net2650 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2716 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_3_575 VPWR VGND sg13g2_fill_1
XFILLER_94_847 VPWR VGND sg13g2_decap_8
XFILLER_59_590 VPWR VGND sg13g2_fill_2
XFILLER_4_1011 VPWR VGND sg13g2_decap_8
XFILLER_93_368 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1263 net2494 net1193 VPWR VGND sg13g2_a22oi_1
XFILLER_47_752 VPWR VGND sg13g2_decap_8
XFILLER_35_903 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2547 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2
+ net2613 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR net650 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_62_733 VPWR VGND sg13g2_fill_1
XFILLER_46_273 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_19_487 VPWR VGND sg13g2_decap_8
XFILLER_62_755 VPWR VGND sg13g2_fill_2
XFILLER_62_744 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\] net627 net2618
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2590 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_43_991 VPWR VGND sg13g2_fill_1
XFILLER_15_671 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_41_clk clknet_5_11__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2628 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y net2755
+ VPWR VGND sg13g2_a22oi_1
XFILLER_61_298 VPWR VGND sg13g2_fill_1
XFILLER_30_641 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2638 i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[364\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net839 net2691 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_30_696 VPWR VGND sg13g2_fill_2
XFILLER_7_870 VPWR VGND sg13g2_fill_1
Xhold837 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\] VPWR
+ VGND net869 sg13g2_dlygate4sd3_1
Xhold804 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] VPWR
+ VGND net836 sg13g2_dlygate4sd3_1
Xhold826 data_pdata\[31\] VPWR VGND net858 sg13g2_dlygate4sd3_1
XFILLER_7_892 VPWR VGND sg13g2_fill_2
XFILLER_6_380 VPWR VGND sg13g2_decap_8
Xhold815 data_pdata\[29\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net847 sg13g2_dlygate4sd3_1
Xhold848 i_snitch.i_snitch_regfile.mem\[52\] VPWR VGND net880 sg13g2_dlygate4sd3_1
Xhold859 i_snitch.i_snitch_regfile.mem\[343\] VPWR VGND net891 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q net3204 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[3\] clknet_leaf_11_clk sg13g2_dfrbpq_2
XFILLER_6_391 VPWR VGND sg13g2_fill_1
Xfanout3290 net3301 net3290 VPWR VGND sg13g2_buf_8
XFILLER_85_836 VPWR VGND sg13g2_decap_8
XFILLER_85_825 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[365\]
+ net3130 i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_65_571 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2889
+ net2653 VPWR VGND sg13g2_nand2_1
XFILLER_52_254 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_32_clk clknet_5_14__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[210\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2792
+ net2675 VPWR VGND sg13g2_nand2_1
XFILLER_4_328 VPWR VGND sg13g2_decap_8
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
XFILLER_106_245 VPWR VGND sg13g2_decap_8
XFILLER_103_963 VPWR VGND sg13g2_decap_8
XFILLER_88_641 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q
+ net3228 VGND VPWR net435 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2777
+ net2660 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_99_clk clknet_5_17__leaf_clk clknet_leaf_99_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2918
+ sg13g2_a221oi_1
XFILLER_48_538 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nor3_2
XFILLER_17_914 VPWR VGND sg13g2_decap_4
XFILLER_84_891 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2388 net1077 net2903 net3039 VPWR VGND sg13g2_a22oi_1
XFILLER_44_755 VPWR VGND sg13g2_decap_4
XFILLER_43_221 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y net2999 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2676
+ net2781 net2273 net2432 VPWR VGND sg13g2_a22oi_1
XFILLER_17_969 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1
+ net777 net618 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_928 VPWR VGND sg13g2_decap_8
XFILLER_106_1011 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_5_12__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2480 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xrsp_state_q_sg13g2_nor2_1_A net914 net2 rsp_state_q_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y VPWR
+ VGND sg13g2_nand2_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_89_1028 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D
+ net3037 net3073 net3147 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B
+ sg13g2_nand4_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y
+ net2815 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ sg13g2_a21oi_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_A1
+ net1363 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2772
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_98_438 VPWR VGND sg13g2_fill_1
XFILLER_98_84 VPWR VGND sg13g2_decap_8
XFILLER_4_884 VPWR VGND sg13g2_decap_4
XFILLER_3_383 VPWR VGND sg13g2_fill_2
XFILLER_94_633 VPWR VGND sg13g2_fill_1
XFILLER_67_869 VPWR VGND sg13g2_fill_2
XFILLER_66_335 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[337\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[414\] clknet_leaf_93_clk sg13g2_dfrbpq_1
XFILLER_82_839 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[203\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[203\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2339 net870 net2679 net2793 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_90_861 VPWR VGND sg13g2_decap_8
XFILLER_62_552 VPWR VGND sg13g2_decap_8
XFILLER_62_574 VPWR VGND sg13g2_fill_1
XFILLER_35_777 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] net3180
+ VPWR VGND sg13g2_nand2b_1
XFILLER_62_596 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2662 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_14_clk clknet_5_6__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B_sg13g2_and2_1_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y
+ net2747 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[15\] net706 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xhold612 i_snitch.i_snitch_regfile.mem\[265\] VPWR VGND net644 sg13g2_dlygate4sd3_1
Xhold601 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net633 sg13g2_dlygate4sd3_1
XFILLER_89_405 VPWR VGND sg13g2_decap_4
Xhold623 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\] VPWR
+ VGND net655 sg13g2_dlygate4sd3_1
Xhold634 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\] VPWR
+ VGND net666 sg13g2_dlygate4sd3_1
Xhold645 data_pdata\[5\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net677 sg13g2_dlygate4sd3_1
XFILLER_104_727 VPWR VGND sg13g2_fill_2
XFILLER_89_438 VPWR VGND sg13g2_fill_2
Xhold667 data_pdata\[4\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net699 sg13g2_dlygate4sd3_1
Xhold678 i_snitch.sb_q\[14\] VPWR VGND net710 sg13g2_dlygate4sd3_1
Xhold656 data_pdata\[3\] VPWR VGND net688 sg13g2_dlygate4sd3_1
Xhold689 data_pdata\[23\] VPWR VGND net721 sg13g2_dlygate4sd3_1
XFILLER_103_259 VPWR VGND sg13g2_decap_8
XFILLER_98_983 VPWR VGND sg13g2_decap_8
XFILLER_58_814 VPWR VGND sg13g2_decap_8
XFILLER_97_482 VPWR VGND sg13g2_decap_8
Xhold1334 rsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1366 sg13g2_dlygate4sd3_1
Xhold1312 rsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1344 sg13g2_dlygate4sd3_1
Xhold1323 i_snitch.inst_addr_o\[18\] VPWR VGND net1355 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1_X
+ VPWR VGND sg13g2_nand2b_1
Xhold1301 i_snitch.i_snitch_regfile.mem\[66\] VPWR VGND net1333 sg13g2_dlygate4sd3_1
XFILLER_100_966 VPWR VGND sg13g2_decap_8
Xhold1356 rsp_data_q\[13\] VPWR VGND net1388 sg13g2_dlygate4sd3_1
Xhold1367 i_req_arb.gen_arbiter.req_d\[1\] VPWR VGND net1399 sg13g2_dlygate4sd3_1
Xhold1345 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\] VPWR
+ VGND net1377 sg13g2_dlygate4sd3_1
Xhold1378 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q VPWR VGND net1410 sg13g2_dlygate4sd3_1
XFILLER_26_722 VPWR VGND sg13g2_decap_8
XFILLER_38_560 VPWR VGND sg13g2_fill_1
XFILLER_81_872 VPWR VGND sg13g2_decap_8
XFILLER_53_585 VPWR VGND sg13g2_fill_1
XFILLER_53_563 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ net3104 VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VGND i_snitch.sb_q\[3\] net2949 sg13g2_o21ai_1
XFILLER_13_416 VPWR VGND sg13g2_fill_2
XFILLER_14_928 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[5\]_sg13g2_dfrbpq_1_Q net3186 VGND VPWR net475 shift_reg_q\[5\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
XFILLER_13_438 VPWR VGND sg13g2_decap_8
XFILLER_13_449 VPWR VGND sg13g2_fill_1
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_B1 VPWR
+ i_snitch.pc_d\[10\] VGND net2305 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_22_972 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2668 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0 net3001 i_snitch.i_snitch_regfile.mem\[130\]
+ i_snitch.i_snitch_regfile.mem\[162\] i_snitch.i_snitch_regfile.mem\[194\] i_snitch.i_snitch_regfile.mem\[226\]
+ net2974 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ net2508 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_49_1001 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[434\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_4_147 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[223\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[223\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2336 net756 net2646 net2790 VPWR VGND sg13g2_a22oi_1
XFILLER_1_832 VPWR VGND sg13g2_decap_8
XFILLER_89_972 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[467\] VGND sg13g2_inv_1
XFILLER_75_110 VPWR VGND sg13g2_fill_2
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_1_1014 VPWR VGND sg13g2_decap_8
XFILLER_17_700 VPWR VGND sg13g2_fill_2
XFILLER_36_519 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[84\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_nand2b_1_A_N_Y
+ net3030 i_snitch.i_snitch_regfile.mem\[84\] VPWR VGND sg13g2_nand2b_1
XFILLER_71_360 VPWR VGND sg13g2_fill_2
XFILLER_17_777 VPWR VGND sg13g2_decap_8
XFILLER_71_382 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VGND net2580 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1293 net2492 net1335 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net673 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2323 net2408 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D net2435
+ sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]
+ net3165 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[114\]
+ net2805 sg13g2_o21ai_1
XFILLER_87_909 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2334
+ sg13g2_o21ai_1
XFILLER_101_708 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[15\]_sg13g2_dfrbpq_1_Q net3232 VGND VPWR rsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[15\] clknet_leaf_35_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_3_clk clknet_5_1__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
XFILLER_95_931 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X
+ net2611 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_or3_1
Xi_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[497\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2365
+ sg13g2_o21ai_1
XFILLER_66_154 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2453 VPWR VGND sg13g2_nand2_1
XFILLER_63_850 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2700 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_90_680 VPWR VGND sg13g2_fill_1
XFILLER_62_393 VPWR VGND sg13g2_fill_1
XFILLER_22_213 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2379
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[454\] clknet_leaf_77_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[302\] net3017 VPWR VGND sg13g2_nand2_1
XFILLER_10_419 VPWR VGND sg13g2_fill_1
XFILLER_22_279 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[243\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[243\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net1023 net2436 net2270 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net701 i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2327 net2485 i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D net2435
+ sg13g2_a221oi_1
Xhold420 i_snitch.i_snitch_regfile.mem\[193\] VPWR VGND net452 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[340\] net2952 VPWR VGND sg13g2_nand2_1
XFILLER_2_607 VPWR VGND sg13g2_decap_8
Xhold442 shift_reg_q\[5\] VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold431 i_snitch.i_snitch_regfile.mem\[129\] VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold453 i_snitch.i_snitch_regfile.mem\[449\] VPWR VGND net485 sg13g2_dlygate4sd3_1
XFILLER_104_524 VPWR VGND sg13g2_fill_2
Xhold464 shift_reg_q\[20\] VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold475 shift_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net507 sg13g2_dlygate4sd3_1
Xhold486 strb_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold497 shift_reg_q\[24\] VPWR VGND net529 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[411\]
+ i_snitch.i_snitch_regfile.mem\[443\] i_snitch.i_snitch_regfile.mem\[475\] i_snitch.i_snitch_regfile.mem\[507\]
+ net3098 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_100_763 VPWR VGND sg13g2_fill_2
XFILLER_86_986 VPWR VGND sg13g2_decap_8
Xhold1142 i_snitch.consec_pc\[0\] VPWR VGND net1174 sg13g2_dlygate4sd3_1
Xhold1120 i_snitch.i_snitch_regfile.mem\[310\] VPWR VGND net1152 sg13g2_dlygate4sd3_1
Xhold1131 i_snitch.i_snitch_regfile.mem\[167\] VPWR VGND net1163 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR net807 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
Xhold1164 i_req_arb.data_i\[42\] VPWR VGND net1196 sg13g2_dlygate4sd3_1
Xhold1175 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\] VPWR
+ VGND net1207 sg13g2_dlygate4sd3_1
Xhold1153 i_snitch.i_snitch_regfile.mem\[426\] VPWR VGND net1185 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_dfrbpq_1_Q_D VGND net2358 net2257
+ sg13g2_o21ai_1
Xhold1197 i_snitch.i_snitch_regfile.mem\[272\] VPWR VGND net1229 sg13g2_dlygate4sd3_1
Xhold1186 i_snitch.i_snitch_regfile.mem\[295\] VPWR VGND net1218 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[72\] VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]
+ net3170 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_81_691 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2414
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_70_22 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y net2695 net2540 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
XFILLER_6_935 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B_Y i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A_X
+ VPWR VGND sg13g2_and4_1
Xi_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_0_161 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2815 VPWR VGND sg13g2_a22oi_1
XFILLER_95_63 VPWR VGND sg13g2_decap_4
XFILLER_77_953 VPWR VGND sg13g2_fill_2
XFILLER_76_452 VPWR VGND sg13g2_decap_8
XFILLER_0_183 VPWR VGND sg13g2_decap_8
XFILLER_92_934 VPWR VGND sg13g2_decap_8
XFILLER_64_636 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[474\] clknet_leaf_116_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1
+ VGND net2610 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C
+ sg13g2_o21ai_1
XFILLER_91_488 VPWR VGND sg13g2_fill_2
XFILLER_91_466 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ net1108 VGND sg13g2_inv_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2760 net2306
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1 net2520 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2323 net1114 net2433 net2284 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ VGND net2600 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2874 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2
+ net2504 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y
+ net114 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_71_190 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B_Y
+ net43 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_728 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_B1 VPWR
+ i_snitch.pc_d\[17\] VGND net2310 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A_Y net3010 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0 net3124 i_snitch.i_snitch_regfile.mem\[137\]
+ i_snitch.i_snitch_regfile.mem\[169\] i_snitch.i_snitch_regfile.mem\[201\] i_snitch.i_snitch_regfile.mem\[233\]
+ net3103 i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[16\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net810 data_pdata\[16\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
XFILLER_99_566 VPWR VGND sg13g2_fill_1
XFILLER_87_728 VPWR VGND sg13g2_decap_4
XFILLER_86_205 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2954 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_68_942 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2366
+ sg13g2_o21ai_1
XFILLER_95_761 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_1 i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_1_Y
+ net2992 i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_nand2b_1_A_N_Y net3021 i_snitch.i_snitch_regfile.mem\[54\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_55_603 VPWR VGND sg13g2_decap_8
XFILLER_83_956 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y
+ VPWR VGND sg13g2_and3_2
XFILLER_50_341 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y
+ net2554 net2602 net2564 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor3_1
XFILLER_23_577 VPWR VGND sg13g2_fill_2
XFILLER_10_238 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_A1 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B
+ VGND VPWR net2533 sg13g2_nor4_2
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0 net3010 i_snitch.i_snitch_regfile.mem\[256\]
+ i_snitch.i_snitch_regfile.mem\[288\] i_snitch.i_snitch_regfile.mem\[320\] i_snitch.i_snitch_regfile.mem\[352\]
+ net2983 i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xfanout3119 net3120 net3119 VPWR VGND sg13g2_buf_8
XFILLER_3_927 VPWR VGND sg13g2_decap_8
Xfanout3108 net3110 net3108 VPWR VGND sg13g2_buf_8
XFILLER_105_833 VPWR VGND sg13g2_decap_8
Xfanout2407 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2407 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[494\] clknet_leaf_83_clk sg13g2_dfrbpq_1
XFILLER_104_343 VPWR VGND sg13g2_decap_8
XFILLER_77_205 VPWR VGND sg13g2_decap_4
Xfanout2429 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y
+ net2429 VPWR VGND sg13g2_buf_8
Xfanout2418 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2418 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_a22oi_1_B2_Y
+ net2323 net670 net2433 net2252 VPWR VGND sg13g2_a22oi_1
XFILLER_49_89 VPWR VGND sg13g2_fill_2
XFILLER_74_901 VPWR VGND sg13g2_fill_2
XFILLER_105_84 VPWR VGND sg13g2_decap_8
XFILLER_58_463 VPWR VGND sg13g2_decap_4
XFILLER_65_66 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[76\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[76\]
+ i_snitch.i_snitch_regfile.mem\[108\] net3133 i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_nor2b_1_Y
+ net3147 net3073 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A
+ VPWR VGND sg13g2_nor2b_1
XFILLER_14_511 VPWR VGND sg13g2_fill_2
XFILLER_26_371 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B net2816
+ i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_81_32 VPWR VGND sg13g2_fill_1
XFILLER_14_533 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1
+ net2867 net2506 i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y VPWR VGND
+ sg13g2_nor3_2
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ VGND net2561 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2554 net2600 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ net2564 sg13g2_a21oi_1
Xi_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X
+ i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q net1331 i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1
+ i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp VPWR VGND
+ sg13g2_a21o_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2700 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_53_8 VPWR VGND sg13g2_fill_2
XFILLER_6_765 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[313\] clknet_leaf_115_clk sg13g2_dfrbpq_1
XFILLER_5_242 VPWR VGND sg13g2_fill_2
XFILLER_5_275 VPWR VGND sg13g2_fill_1
XFILLER_69_717 VPWR VGND sg13g2_decap_8
XFILLER_69_706 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2411 net1072 net2900 net2870 VPWR VGND sg13g2_a22oi_1
Xfanout2930 net2932 net2930 VPWR VGND sg13g2_buf_8
XFILLER_96_547 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B VPWR
+ VGND sg13g2_nor3_1
XFILLER_69_739 VPWR VGND sg13g2_fill_1
Xfanout2952 net2953 net2952 VPWR VGND sg13g2_buf_8
Xfanout2941 net2946 net2941 VPWR VGND sg13g2_buf_8
XFILLER_2_971 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_nor3_1_A net1279 net2764 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xfanout2963 net2966 net2963 VPWR VGND sg13g2_buf_8
Xfanout2996 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ net2996 VPWR VGND sg13g2_buf_8
Xfanout2985 net2986 net2985 VPWR VGND sg13g2_buf_8
Xfanout2974 net2976 net2974 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[419\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[419\]
+ net3006 i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_a21oi_1_A1_Y net2979 sg13g2_a21oi_1
XFILLER_77_794 VPWR VGND sg13g2_fill_1
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_64_400 VPWR VGND sg13g2_fill_1
XFILLER_37_614 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_A1
+ net1401 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2357
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
XFILLER_64_466 VPWR VGND sg13g2_decap_8
XFILLER_52_606 VPWR VGND sg13g2_fill_1
XFILLER_80_959 VPWR VGND sg13g2_decap_8
XFILLER_52_639 VPWR VGND sg13g2_decap_8
XFILLER_51_116 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[309\]
+ net2810 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[385\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net495 net2389 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0_X net2954 i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_mux4_1_A0_X sg13g2_a221oi_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2593 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1_sg13g2_nor4_1_Y
+ net3079 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D
+ net96 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor4_1
Xshift_reg_q\[9\]_sg13g2_a22oi_1_A1 shift_reg_q\[9\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_mux2_1_A1_1_X
+ net3054 net3044 shift_reg_q\[9\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_341 VPWR VGND sg13g2_fill_1
XFILLER_0_919 VPWR VGND sg13g2_decap_8
XFILLER_102_814 VPWR VGND sg13g2_decap_8
XFILLER_87_536 VPWR VGND sg13g2_fill_1
XFILLER_101_357 VPWR VGND sg13g2_decap_8
XFILLER_19_15 VPWR VGND sg13g2_fill_2
XFILLER_67_260 VPWR VGND sg13g2_fill_1
XFILLER_83_731 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_nand3b_1_B_Y
+ sg13g2_a221oi_1
XFILLER_83_786 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net801 net2651 net2863 VPWR VGND sg13g2_a22oi_1
XFILLER_55_488 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[291\] VGND sg13g2_inv_1
XFILLER_36_680 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q
+ net3234 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[500\]_sg13g2_o21ai_1_A1 net2965 VPWR i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[500\] net2806 sg13g2_o21ai_1
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[333\] clknet_leaf_85_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2448 net2255 net2409 net1250 VPWR VGND sg13g2_a22oi_1
XFILLER_51_79 VPWR VGND sg13g2_fill_1
XFILLER_7_518 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B
+ sg13g2_o21ai_1
XFILLER_104_140 VPWR VGND sg13g2_decap_8
XFILLER_78_503 VPWR VGND sg13g2_fill_2
XFILLER_3_779 VPWR VGND sg13g2_decap_4
Xfanout2237 net2237 net2238 VPWR VGND sg13g2_buf_16
Xfanout2248 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y
+ net2248 VPWR VGND sg13g2_buf_8
Xfanout2259 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2259 VPWR VGND sg13g2_buf_8
Xshift_reg_q\[21\]_sg13g2_a22oi_1_A1 shift_reg_q\[21\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_1_X
+ net3053 net3043 shift_reg_q\[21\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_58_260 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_o21ai_1_A2
+ net3054 VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ VGND net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]
+ sg13g2_o21ai_1
XFILLER_76_98 VPWR VGND sg13g2_fill_2
XFILLER_74_720 VPWR VGND sg13g2_decap_8
XFILLER_58_271 VPWR VGND sg13g2_fill_1
XFILLER_19_647 VPWR VGND sg13g2_fill_1
XFILLER_20_1018 VPWR VGND sg13g2_decap_8
XFILLER_74_753 VPWR VGND sg13g2_decap_8
XFILLER_19_669 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2958
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2963
+ i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
XFILLER_15_831 VPWR VGND sg13g2_fill_2
XFILLER_33_116 VPWR VGND sg13g2_fill_1
XFILLER_15_842 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_A1
+ net2309 i_snitch.pc_d\[23\] i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2632 VPWR i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2636 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_97_845 VPWR VGND sg13g2_decap_8
XFILLER_97_812 VPWR VGND sg13g2_fill_1
XFILLER_69_525 VPWR VGND sg13g2_decap_8
Xfanout2760 net2763 net2760 VPWR VGND sg13g2_buf_8
XFILLER_69_547 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xfanout2771 net2772 net2771 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2597 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X net3
+ i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S VPWR VGND sg13g2_mux2_1
XFILLER_84_528 VPWR VGND sg13g2_fill_2
XFILLER_84_506 VPWR VGND sg13g2_fill_1
XFILLER_56_208 VPWR VGND sg13g2_fill_2
Xfanout2782 net2783 net2782 VPWR VGND sg13g2_buf_8
Xfanout2793 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1_X
+ net2793 VPWR VGND sg13g2_buf_8
XFILLER_84_539 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[353\] clknet_leaf_76_clk sg13g2_dfrbpq_1
Xdata_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1 data_pdata\[15\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y
+ data_pdata\[15\]_sg13g2_nand2b_1_B_Y data_pdata\[23\]_sg13g2_a21oi_1_A2_Y data_pdata\[31\]_sg13g2_nand2b_1_B_Y
+ net3152 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net1116 net2688 net2889 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2604 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_25_617 VPWR VGND sg13g2_decap_8
XFILLER_25_628 VPWR VGND sg13g2_fill_1
XFILLER_80_756 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C
+ net2923 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_and3_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[62\]
+ net2986 sg13g2_o21ai_1
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ VGND VPWR net39 sg13g2_nor4_2
XFILLER_20_333 VPWR VGND sg13g2_fill_1
XFILLER_32_182 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2733 shift_reg_q\[23\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[19\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[19\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_20_399 VPWR VGND sg13g2_decap_8
XFILLER_21_27 VPWR VGND sg13g2_fill_2
XFILLER_106_427 VPWR VGND sg13g2_decap_8
Xdata_pdata\[2\]_sg13g2_mux2_1_A1 rsp_data_q\[2\] net686 net3048 data_pdata\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_99_171 VPWR VGND sg13g2_decap_8
XFILLER_99_160 VPWR VGND sg13g2_fill_2
XFILLER_0_716 VPWR VGND sg13g2_decap_8
XFILLER_102_655 VPWR VGND sg13g2_decap_8
XFILLER_87_344 VPWR VGND sg13g2_fill_2
XFILLER_87_333 VPWR VGND sg13g2_fill_2
XFILLER_101_154 VPWR VGND sg13g2_decap_8
XFILLER_88_889 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[13\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.pc_d\[13\]
+ i_snitch.inst_addr_o\[13\] clknet_leaf_53_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[328\] VGND sg13g2_inv_1
XFILLER_83_594 VPWR VGND sg13g2_decap_8
XFILLER_16_628 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2605 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_102_63 VPWR VGND sg13g2_decap_8
XFILLER_71_767 VPWR VGND sg13g2_fill_2
XFILLER_71_778 VPWR VGND sg13g2_fill_2
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_7_18 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[478\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net935 net2461 net2244 VPWR VGND sg13g2_a22oi_1
XFILLER_7_348 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q
+ net3240 VGND VPWR net961 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[373\] clknet_leaf_114_clk sg13g2_dfrbpq_1
XFILLER_106_983 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ net2584 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_78_311 VPWR VGND sg13g2_decap_8
XFILLER_78_344 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2825
+ sg13g2_a221oi_1
XFILLER_93_303 VPWR VGND sg13g2_fill_1
XFILLER_78_388 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[479\]
+ net2949 i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_a21o_1_A1_X
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y
+ net46 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B
+ VPWR VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y
+ sg13g2_nand3b_1
XFILLER_66_539 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2845
+ sg13g2_a221oi_1
XFILLER_35_926 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[369\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[369\] net2807 sg13g2_o21ai_1
XFILLER_43_981 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[508\] clknet_leaf_95_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold805 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net837 sg13g2_dlygate4sd3_1
Xhold827 data_pdata\[31\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net859 sg13g2_dlygate4sd3_1
Xhold816 i_snitch.i_snitch_regfile.mem\[363\] VPWR VGND net848 sg13g2_dlygate4sd3_1
XFILLER_6_370 VPWR VGND sg13g2_fill_2
Xhold849 i_snitch.i_snitch_regfile.mem\[470\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold838 i_snitch.i_snitch_regfile.mem\[203\] VPWR VGND net870 sg13g2_dlygate4sd3_1
XFILLER_97_653 VPWR VGND sg13g2_fill_1
XFILLER_97_631 VPWR VGND sg13g2_decap_8
Xfanout3291 net3300 net3291 VPWR VGND sg13g2_buf_8
Xfanout3280 net3281 net3280 VPWR VGND sg13g2_buf_8
Xfanout2590 net2591 net2590 VPWR VGND sg13g2_buf_8
XFILLER_93_881 VPWR VGND sg13g2_decap_8
XFILLER_53_712 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[498\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2458 net2273 net2369 net1261 VPWR VGND sg13g2_a22oi_1
XFILLER_37_263 VPWR VGND sg13g2_decap_8
XFILLER_38_797 VPWR VGND sg13g2_decap_4
XFILLER_80_542 VPWR VGND sg13g2_fill_1
XFILLER_52_222 VPWR VGND sg13g2_decap_8
XFILLER_16_38 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[393\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_21_620 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q
+ net3184 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_34_992 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_nand2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y net2817
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C i_snitch.inst_addr_o\[21\]
+ net2308 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_B1
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[182\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net1045 net2651 net2775 VPWR VGND sg13g2_a22oi_1
XFILLER_10_1006 VPWR VGND sg13g2_decap_8
XFILLER_106_224 VPWR VGND sg13g2_decap_8
XFILLER_103_942 VPWR VGND sg13g2_decap_8
XFILLER_87_163 VPWR VGND sg13g2_fill_2
XFILLER_57_45 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_29_731 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[317\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2431 net2251 net2317 net1211 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ net2582 VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ VGND net2597 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ sg13g2_o21ai_1
XFILLER_84_870 VPWR VGND sg13g2_decap_8
XFILLER_56_561 VPWR VGND sg13g2_fill_1
XFILLER_16_403 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q net3323 VGND VPWR i_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[212\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_43_277 VPWR VGND sg13g2_fill_2
Xstrb_reg_q\[0\]_sg13g2_a22oi_1_A1 strb_out_sg13g2_inv_1_Y_A strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B2 cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 strb_reg_q\[0\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2721 i_snitch.inst_addr_o\[25\] sg13g2_a21oi_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_B1
+ VGND VPWR i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A_Y
+ target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q_D
+ net125 sg13g2_a21oi_1
XFILLER_24_480 VPWR VGND sg13g2_decap_4
XFILLER_12_653 VPWR VGND sg13g2_fill_2
XFILLER_89_1007 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[318\]
+ net3015 i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_a21oi_1_A1_Y net2986 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B
+ net95 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ net2719 i_req_arb.data_i\[37\] VPWR VGND sg13g2_a22oi_1
XFILLER_106_780 VPWR VGND sg13g2_decap_8
XFILLER_98_63 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2959
+ i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2965
+ i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
XFILLER_3_351 VPWR VGND sg13g2_decap_4
Xstrb_reg_q\[1\]_sg13g2_a21oi_1_A1 VGND VPWR strb_reg_q\[1\] net3044 strb_reg_q\[1\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B2 sg13g2_a21oi_1
Xdata_pdata\[9\]_sg13g2_mux2_1_A1 rsp_data_q\[9\] net889 net3048 data_pdata\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_94_645 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[10\] net1003 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_67_859 VPWR VGND sg13g2_fill_1
XFILLER_67_848 VPWR VGND sg13g2_decap_8
XFILLER_94_656 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xtarget_sel_q_sg13g2_nor2_1_A net1026 target_sel_q_sg13g2_nor2_1_A_B target_sel_q_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_93_177 VPWR VGND sg13g2_fill_2
XFILLER_75_892 VPWR VGND sg13g2_decap_8
Xcnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2_1_Y cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A
+ net1 cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 VPWR VGND sg13g2_nand2_2
XFILLER_90_840 VPWR VGND sg13g2_decap_8
XFILLER_50_704 VPWR VGND sg13g2_decap_4
XFILLER_72_1000 VPWR VGND sg13g2_fill_2
XFILLER_16_992 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_962 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_mux2_1_A0_X net3108 net2827 i_snitch.i_snitch_regfile.mem\[50\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_33_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1076 net2456 net2273 VPWR VGND sg13g2_a22oi_1
Xhold602 i_snitch.i_snitch_regfile.mem\[264\] VPWR VGND net634 sg13g2_dlygate4sd3_1
Xhold635 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\] VPWR
+ VGND net667 sg13g2_dlygate4sd3_1
Xhold613 i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND net645 sg13g2_dlygate4sd3_1
Xhold624 i_snitch.i_snitch_regfile.mem\[335\] VPWR VGND net656 sg13g2_dlygate4sd3_1
Xhold679 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net711 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2404 net723 net2663 net2797 VPWR VGND sg13g2_a22oi_1
Xhold668 i_snitch.i_snitch_regfile.mem\[281\] VPWR VGND net700 sg13g2_dlygate4sd3_1
Xhold646 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_inv_1_A_Y VPWR VGND net678 sg13g2_dlygate4sd3_1
Xhold657 data_pdata\[3\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net689 sg13g2_dlygate4sd3_1
XFILLER_103_238 VPWR VGND sg13g2_decap_8
XFILLER_98_962 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1 net3022 i_snitch.i_snitch_regfile.mem\[151\]
+ i_snitch.i_snitch_regfile.mem\[183\] i_snitch.i_snitch_regfile.mem\[215\] i_snitch.i_snitch_regfile.mem\[247\]
+ net2993 i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2868
+ net2656 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2442 net2773 i_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
XFILLER_100_945 VPWR VGND sg13g2_decap_8
Xhold1313 rsp_data_q\[27\] VPWR VGND net1345 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[232\] clknet_leaf_73_clk sg13g2_dfrbpq_1
Xhold1324 i_snitch.i_snitch_regfile.mem\[423\] VPWR VGND net1356 sg13g2_dlygate4sd3_1
Xhold1302 i_snitch.i_snitch_regfile.mem\[354\] VPWR VGND net1334 sg13g2_dlygate4sd3_1
XFILLER_85_667 VPWR VGND sg13g2_fill_2
XFILLER_85_656 VPWR VGND sg13g2_fill_2
Xhold1368 i_snitch.inst_addr_o\[12\] VPWR VGND net1400 sg13g2_dlygate4sd3_1
Xhold1346 i_req_arb.data_i\[37\] VPWR VGND net1378 sg13g2_dlygate4sd3_1
Xhold1357 i_snitch.gpr_waddr\[7\] VPWR VGND net1389 sg13g2_dlygate4sd3_1
Xhold1335 i_snitch.gpr_waddr\[6\] VPWR VGND net1367 sg13g2_dlygate4sd3_1
XFILLER_72_328 VPWR VGND sg13g2_decap_8
XFILLER_81_851 VPWR VGND sg13g2_decap_8
XFILLER_65_391 VPWR VGND sg13g2_fill_2
XFILLER_25_244 VPWR VGND sg13g2_decap_8
XFILLER_80_394 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\] net589 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xtarget_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y req_data_valid_sg13g2_o21ai_1_Y_B1
+ target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B target_sel_q_sg13g2_nor2_1_A_B
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_nand2_1_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_nand2_1_A_Y
+ net428 net2616 VPWR VGND sg13g2_nand2_1
XFILLER_5_649 VPWR VGND sg13g2_fill_1
XFILLER_4_126 VPWR VGND sg13g2_decap_8
XFILLER_1_811 VPWR VGND sg13g2_decap_8
XFILLER_89_951 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_C1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B_Y
+ sg13g2_a21oi_1
XFILLER_88_450 VPWR VGND sg13g2_fill_1
XFILLER_0_332 VPWR VGND sg13g2_fill_2
XFILLER_1_888 VPWR VGND sg13g2_decap_8
XFILLER_88_472 VPWR VGND sg13g2_decap_4
XFILLER_76_634 VPWR VGND sg13g2_fill_1
XFILLER_48_314 VPWR VGND sg13g2_fill_1
XFILLER_0_365 VPWR VGND sg13g2_decap_8
XFILLER_48_369 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2745 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_17_723 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2713 i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_95_1022 VPWR VGND sg13g2_decap_8
XFILLER_75_199 VPWR VGND sg13g2_fill_2
XFILLER_57_892 VPWR VGND sg13g2_fill_1
XFILLER_16_222 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net1103 net2900 net2786 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2700 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1_Y
+ sg13g2_a21oi_1
XFILLER_31_236 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2885
+ net2657 VPWR VGND sg13g2_nand2_1
XFILLER_12_494 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] net630 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1 net3000 i_snitch.i_snitch_regfile.mem\[153\]
+ i_snitch.i_snitch_regfile.mem\[185\] i_snitch.i_snitch_regfile.mem\[217\] i_snitch.i_snitch_regfile.mem\[249\]
+ net2973 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_9_999 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1_sg13g2_and2_1_X
+ net3144 net3142 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[252\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[71\]
+ net2841 i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
XFILLER_99_726 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1 VPWR VGND net3109 net2822
+ i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[46\]
+ i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1_Y net2830 sg13g2_a221oi_1
XFILLER_4_682 VPWR VGND sg13g2_fill_2
XFILLER_95_910 VPWR VGND sg13g2_decap_8
XFILLER_79_461 VPWR VGND sg13g2_fill_2
XFILLER_100_219 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[358\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[358\]
+ net124 i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
XFILLER_39_325 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2545 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2611 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[202\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_987 VPWR VGND sg13g2_decap_8
XFILLER_94_464 VPWR VGND sg13g2_decap_4
XFILLER_81_114 VPWR VGND sg13g2_fill_2
XFILLER_66_188 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_63_884 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1 VPWR VGND i_snitch.inst_addr_o\[27\]
+ i_snitch.pc_d\[18\]_sg13g2_mux2_1_A1_X net56 i_snitch.inst_addr_o\[22\] i_snitch.pc_d\[18\]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_inv_1_A_Y sg13g2_a221oi_1
XFILLER_63_895 VPWR VGND sg13g2_decap_8
XFILLER_50_512 VPWR VGND sg13g2_decap_4
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
XFILLER_23_759 VPWR VGND sg13g2_fill_2
XFILLER_13_39 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1343 net3065 rsp_data_q\[5\] VPWR VGND sg13g2_a22oi_1
XFILLER_31_792 VPWR VGND sg13g2_fill_1
Xhold410 strb_reg_q\[6\] VPWR VGND net442 sg13g2_dlygate4sd3_1
Xhold454 shift_reg_q\[14\] VPWR VGND net486 sg13g2_dlygate4sd3_1
Xhold421 i_snitch.i_snitch_regfile.mem\[510\] VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold443 shift_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold432 i_snitch.i_snitch_regfile.mem\[161\] VPWR VGND net464 sg13g2_dlygate4sd3_1
XFILLER_104_547 VPWR VGND sg13g2_fill_1
XFILLER_89_214 VPWR VGND sg13g2_fill_1
Xhold465 shift_reg_q\[20\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net497 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q_D VGND net2259 net2386
+ sg13g2_o21ai_1
Xhold476 shift_reg_q\[18\] VPWR VGND net508 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_dfrbpq_1_Q
+ net3191 VGND VPWR net588 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
Xhold487 shift_reg_q\[11\] VPWR VGND net519 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
Xhold498 shift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net530 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net1110 net2451 net2255 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2b_1_Y
+ req_data_valid_sg13g2_o21ai_1_Y_B1 target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_nor2b_1
XFILLER_86_965 VPWR VGND sg13g2_decap_8
XFILLER_85_453 VPWR VGND sg13g2_decap_8
Xhold1121 rsp_data_q\[15\] VPWR VGND net1153 sg13g2_dlygate4sd3_1
XFILLER_58_667 VPWR VGND sg13g2_decap_4
Xhold1110 i_snitch.i_snitch_regfile.mem\[143\] VPWR VGND net1142 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2771
+ net2659 VPWR VGND sg13g2_nand2_1
Xhold1132 i_snitch.i_snitch_regfile.mem\[402\] VPWR VGND net1164 sg13g2_dlygate4sd3_1
XFILLER_79_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1 VPWR VGND i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_C1 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y
+ i_snitch.inst_addr_o\[18\] i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_Y net2724
+ sg13g2_a221oi_1
XFILLER_73_604 VPWR VGND sg13g2_decap_8
Xhold1165 i_snitch.inst_addr_o\[25\] VPWR VGND net1197 sg13g2_dlygate4sd3_1
Xhold1143 i_snitch.i_snitch_regfile.mem\[181\] VPWR VGND net1175 sg13g2_dlygate4sd3_1
Xhold1154 i_snitch.i_snitch_regfile.mem\[441\] VPWR VGND net1186 sg13g2_dlygate4sd3_1
Xhold1176 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] VPWR
+ VGND net1208 sg13g2_dlygate4sd3_1
Xhold1198 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] VPWR
+ VGND net1230 sg13g2_dlygate4sd3_1
XFILLER_45_339 VPWR VGND sg13g2_fill_1
XFILLER_45_328 VPWR VGND sg13g2_decap_8
Xhold1187 i_snitch.i_snitch_regfile.mem\[67\] VPWR VGND net1219 sg13g2_dlygate4sd3_1
XFILLER_81_670 VPWR VGND sg13g2_fill_1
XFILLER_53_372 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1 net2999 i_snitch.i_snitch_regfile.mem\[155\]
+ i_snitch.i_snitch_regfile.mem\[187\] i_snitch.i_snitch_regfile.mem\[219\] i_snitch.i_snitch_regfile.mem\[251\]
+ net2973 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_13_258 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[272\] clknet_leaf_87_clk sg13g2_dfrbpq_1
XFILLER_41_545 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_or3_1_X
+ net96 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B
+ VPWR VGND sg13g2_or3_1
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1 VPWR VGND net3108 net2822
+ i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[48\]
+ i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1_Y net2827 sg13g2_a221oi_1
XFILLER_22_781 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2731 shift_reg_q\[11\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[7\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[7\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_103_1026 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1336 net2492 net1287 VPWR VGND sg13g2_a22oi_1
XFILLER_6_903 VPWR VGND sg13g2_fill_2
XFILLER_10_932 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2703 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A
+ net3081 net3075 VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ net2626 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[378\]
+ net3116 i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_102_0 VPWR VGND sg13g2_decap_8
XFILLER_79_21 VPWR VGND sg13g2_fill_1
XFILLER_5_479 VPWR VGND sg13g2_fill_2
XFILLER_79_65 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[13\]_sg13g2_nor2_1_A net476 net2728 shift_reg_q\[13\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[300\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_dfrbpq_1_Q_D VGND net2393 net310
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_B_sg13g2_inv_1_Y VPWR i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_B
+ i_snitch.i_snitch_lsu.metadata_q\[1\] VGND sg13g2_inv_1
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_B1
+ net668 net2785 VPWR VGND sg13g2_nand2b_1
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2783 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2
+ net2506 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_2
XFILLER_62_1021 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[268\]_sg13g2_o21ai_1_A1 net2937 VPWR i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[268\] net2814 sg13g2_o21ai_1
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_1_685 VPWR VGND sg13g2_decap_8
XFILLER_95_42 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[407\] clknet_leaf_67_clk sg13g2_dfrbpq_1
XFILLER_0_195 VPWR VGND sg13g2_decap_8
XFILLER_92_913 VPWR VGND sg13g2_decap_8
XFILLER_77_998 VPWR VGND sg13g2_decap_8
XFILLER_91_434 VPWR VGND sg13g2_decap_8
XFILLER_29_391 VPWR VGND sg13g2_decap_4
XFILLER_63_147 VPWR VGND sg13g2_fill_1
XFILLER_45_862 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[282\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2697 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_32_556 VPWR VGND sg13g2_decap_8
XFILLER_32_567 VPWR VGND sg13g2_fill_1
XFILLER_60_887 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D_sg13g2_and4_1_X
+ net3035 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D
+ VPWR VGND sg13g2_and4_1
XFILLER_9_741 VPWR VGND sg13g2_fill_2
Xcnt_q\[1\]_sg13g2_dfrbpq_1_Q net3184 VGND VPWR cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D cnt_q\[1\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ net2631 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y
+ net2576 net2564 net59 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_Y
+ VPWR VGND i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A
+ sg13g2_nand4_1
XFILLER_5_991 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2435 VPWR VGND sg13g2_nand2_1
XFILLER_99_556 VPWR VGND sg13g2_fill_1
XFILLER_5_95 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2389 net850 net2689 net3040 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2456 VPWR VGND sg13g2_nand2_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y VPWR
+ VGND sg13g2_nor3_2
XFILLER_95_740 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2627 net2758 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_a22oi_1
XFILLER_68_965 VPWR VGND sg13g2_fill_2
XFILLER_67_420 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1 net3012 i_snitch.i_snitch_regfile.mem\[157\]
+ i_snitch.i_snitch_regfile.mem\[189\] i_snitch.i_snitch_regfile.mem\[221\] i_snitch.i_snitch_regfile.mem\[253\]
+ net2985 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[259\]_sg13g2_nor3_1_A net1359 net2892 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_83_935 VPWR VGND sg13g2_decap_8
XFILLER_68_987 VPWR VGND sg13g2_fill_2
XFILLER_27_306 VPWR VGND sg13g2_decap_4
XFILLER_28_829 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[292\] clknet_leaf_109_clk sg13g2_dfrbpq_1
XFILLER_94_283 VPWR VGND sg13g2_fill_2
XFILLER_82_467 VPWR VGND sg13g2_fill_1
XFILLER_36_851 VPWR VGND sg13g2_fill_2
XFILLER_36_862 VPWR VGND sg13g2_decap_8
XFILLER_36_873 VPWR VGND sg13g2_fill_2
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[288\]_sg13g2_o21ai_1_A1 net2939 VPWR i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[288\] net2811 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[427\] clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_40_37 VPWR VGND sg13g2_fill_1
XFILLER_105_812 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y
+ net2574 VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ VGND net2581 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
Xshift_reg_q\[26\]_sg13g2_nor2_1_A net550 net2734 shift_reg_q\[26\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_906 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2742
+ net2649 VPWR VGND sg13g2_nand2_1
Xfanout3109 net3110 net3109 VPWR VGND sg13g2_buf_8
XFILLER_104_322 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[216\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[216\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net808 net2666 net2791 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q_D VGND net2521 net2328
+ sg13g2_o21ai_1
XFILLER_6_7 VPWR VGND sg13g2_decap_8
Xfanout2408 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2408 VPWR VGND sg13g2_buf_8
XFILLER_105_889 VPWR VGND sg13g2_decap_8
Xfanout2419 net2420 net2419 VPWR VGND sg13g2_buf_2
XFILLER_46_1027 VPWR VGND sg13g2_fill_2
XFILLER_46_1016 VPWR VGND sg13g2_decap_8
XFILLER_104_399 VPWR VGND sg13g2_decap_8
XFILLER_59_943 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[111\] clknet_leaf_63_clk sg13g2_dfrbpq_1
XFILLER_105_63 VPWR VGND sg13g2_decap_8
XFILLER_100_594 VPWR VGND sg13g2_fill_1
XFILLER_46_648 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0 net3130 i_snitch.i_snitch_regfile.mem\[141\]
+ i_snitch.i_snitch_regfile.mem\[173\] i_snitch.i_snitch_regfile.mem\[205\] i_snitch.i_snitch_regfile.mem\[237\]
+ net3108 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_xor2_1
XFILLER_92_1025 VPWR VGND sg13g2_decap_4
XFILLER_61_629 VPWR VGND sg13g2_fill_1
XFILLER_60_106 VPWR VGND sg13g2_fill_1
XFILLER_81_22 VPWR VGND sg13g2_fill_1
XFILLER_14_545 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2538 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ net2572 sg13g2_a21oi_2
Xrsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1226 net3067 rsp_data_q\[14\] VPWR VGND sg13g2_a22oi_1
Xshift_reg_q\[10\]_sg13g2_dfrbpq_1_Q net3198 VGND VPWR net469 shift_reg_q\[10\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_42_887 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y net2512
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_14_71 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2
+ VGND VPWR net3165 net606 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1 net3009 i_snitch.i_snitch_regfile.mem\[159\]
+ i_snitch.i_snitch_regfile.mem\[191\] i_snitch.i_snitch_regfile.mem\[223\] i_snitch.i_snitch_regfile.mem\[255\]
+ net2982 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_2_950 VPWR VGND sg13g2_decap_8
Xfanout2920 net2920 net2921 VPWR VGND sg13g2_buf_16
XFILLER_68_228 VPWR VGND sg13g2_fill_2
Xfanout2953 net111 net2953 VPWR VGND sg13g2_buf_8
Xfanout2931 net2932 net2931 VPWR VGND sg13g2_buf_8
XFILLER_1_460 VPWR VGND sg13g2_decap_8
Xfanout2942 net2945 net2942 VPWR VGND sg13g2_buf_8
Xfanout2964 net2966 net2964 VPWR VGND sg13g2_buf_8
XFILLER_77_751 VPWR VGND sg13g2_fill_1
Xfanout2997 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2997 VPWR VGND sg13g2_buf_8
XFILLER_49_431 VPWR VGND sg13g2_decap_4
Xfanout2975 net2976 net2975 VPWR VGND sg13g2_buf_1
Xfanout2986 net2995 net2986 VPWR VGND sg13g2_buf_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_77_762 VPWR VGND sg13g2_fill_1
XFILLER_49_475 VPWR VGND sg13g2_decap_8
XFILLER_92_721 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_49_497 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0 net3122 i_snitch.i_snitch_regfile.mem\[260\]
+ i_snitch.i_snitch_regfile.mem\[292\] i_snitch.i_snitch_regfile.mem\[324\] i_snitch.i_snitch_regfile.mem\[356\]
+ net3104 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2554 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_36_169 VPWR VGND sg13g2_fill_1
XFILLER_80_938 VPWR VGND sg13g2_decap_8
XFILLER_51_128 VPWR VGND sg13g2_decap_8
XFILLER_51_106 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ net92 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y
+ sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q net3305 VGND VPWR i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[447\] clknet_leaf_53_clk sg13g2_dfrbpq_2
XFILLER_51_139 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ net33 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2
+ VPWR VGND sg13g2_nor3_1
XFILLER_33_898 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[236\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[236\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net1056 net2692 net2875 VPWR VGND sg13g2_a22oi_1
XFILLER_60_695 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[80\]
+ i_snitch.i_snitch_regfile.mem\[112\] net3131 i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2891 net2912 i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_10_18 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2 net2832
+ VPWR i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[131\] clknet_leaf_108_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2
+ net2507 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_105_119 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1
+ VGND VPWR net2744 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2392
+ sg13g2_o21ai_1
XFILLER_99_386 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net2557 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
XFILLER_101_336 VPWR VGND sg13g2_decap_8
XFILLER_95_592 VPWR VGND sg13g2_decap_4
XFILLER_83_765 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2761 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_43_607 VPWR VGND sg13g2_fill_1
XFILLER_35_15 VPWR VGND sg13g2_fill_1
XFILLER_55_478 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y net3000 sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2481 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_51_651 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2713 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[28\]_sg13g2_dfrbpq_1_Q net3243 VGND VPWR rsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[28\] clknet_leaf_33_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A_Y net2953 i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2945 sg13g2_a21oi_1
XFILLER_105_620 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_nor2_1_A
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A net2626
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_C1
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_714 VPWR VGND sg13g2_decap_8
XFILLER_3_758 VPWR VGND sg13g2_decap_8
XFILLER_2_246 VPWR VGND sg13g2_fill_2
Xfanout2238 net2238 net2241 VPWR VGND sg13g2_buf_16
Xfanout2249 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y
+ net2249 VPWR VGND sg13g2_buf_8
XFILLER_104_196 VPWR VGND sg13g2_decap_8
XFILLER_78_548 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2458
+ net2514 net2902 net2857 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B
+ net2566 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[467\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[432\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net438 net2381 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[162\]_sg13g2_nor3_1_A net1282 net2772 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[162\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_100_380 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_92_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2323 net865 net2904 net2892 VPWR VGND sg13g2_a22oi_1
XFILLER_74_798 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[151\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_26_180 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y
+ net2612 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B
+ VPWR VGND sg13g2_nand2_2
XFILLER_70_971 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[470\] net2952 VPWR VGND sg13g2_nand2_1
XFILLER_25_92 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1
+ VPWR VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_C1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X
+ sg13g2_a221oi_1
XFILLER_97_824 VPWR VGND sg13g2_decap_8
Xfanout2750 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2750 VPWR VGND sg13g2_buf_8
Xfanout2761 net2763 net2761 VPWR VGND sg13g2_buf_8
XFILLER_2_791 VPWR VGND sg13g2_fill_1
Xfanout2772 net2773 net2772 VPWR VGND sg13g2_buf_8
Xfanout2794 net2799 net2794 VPWR VGND sg13g2_buf_8
Xfanout2783 net2784 net2783 VPWR VGND sg13g2_buf_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_65_765 VPWR VGND sg13g2_fill_2
XFILLER_64_242 VPWR VGND sg13g2_decap_4
XFILLER_53_905 VPWR VGND sg13g2_fill_2
XFILLER_49_294 VPWR VGND sg13g2_decap_8
XFILLER_38_979 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2695 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_80_724 VPWR VGND sg13g2_fill_2
XFILLER_52_426 VPWR VGND sg13g2_fill_2
XFILLER_52_415 VPWR VGND sg13g2_decap_8
XFILLER_24_117 VPWR VGND sg13g2_fill_1
XFILLER_75_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0 net3138 i_snitch.i_snitch_regfile.mem\[148\]
+ i_snitch.i_snitch_regfile.mem\[180\] i_snitch.i_snitch_regfile.mem\[212\] i_snitch.i_snitch_regfile.mem\[244\]
+ net3111 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_52_437 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ VGND net2709 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B net2301 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
XFILLER_61_982 VPWR VGND sg13g2_decap_4
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
XFILLER_106_406 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_Y
+ net3141 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_1 i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_1_Y
+ net2977 i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_nand2b_1_A_N_Y net3004 i_snitch.i_snitch_regfile.mem\[59\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[487\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[276\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2325 net785 net2672 net2893 VPWR VGND sg13g2_a22oi_1
XFILLER_99_194 VPWR VGND sg13g2_fill_1
XFILLER_88_868 VPWR VGND sg13g2_decap_8
XFILLER_101_133 VPWR VGND sg13g2_decap_8
XFILLER_75_507 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[171\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_56_754 VPWR VGND sg13g2_decap_4
XFILLER_55_220 VPWR VGND sg13g2_decap_4
XFILLER_46_36 VPWR VGND sg13g2_fill_2
XFILLER_29_968 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND net2580 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_46_69 VPWR VGND sg13g2_fill_1
XFILLER_102_42 VPWR VGND sg13g2_decap_8
XFILLER_70_245 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0 net3135 i_snitch.i_snitch_regfile.mem\[267\]
+ i_snitch.i_snitch_regfile.mem\[299\] i_snitch.i_snitch_regfile.mem\[331\] i_snitch.i_snitch_regfile.mem\[363\]
+ net3112 i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[29\]_sg13g2_dfrbpq_1_Q net3191 VGND VPWR net847 data_pdata\[29\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
XFILLER_8_817 VPWR VGND sg13g2_fill_1
XFILLER_7_305 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1299 net3066 rsp_data_q\[3\] VPWR VGND sg13g2_a22oi_1
XFILLER_7_338 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2933 i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[306\] clknet_leaf_93_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[87\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[87\]
+ i_snitch.i_snitch_regfile.mem\[119\] net3138 i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_106_962 VPWR VGND sg13g2_decap_8
XFILLER_11_72 VPWR VGND sg13g2_fill_1
XFILLER_79_802 VPWR VGND sg13g2_fill_2
XFILLER_78_367 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_59_592 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1_X net2964 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2706 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_19_467 VPWR VGND sg13g2_fill_2
XFILLER_74_595 VPWR VGND sg13g2_decap_8
XFILLER_62_757 VPWR VGND sg13g2_fill_1
XFILLER_34_426 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0 net3001 i_snitch.i_snitch_regfile.mem\[386\]
+ i_snitch.i_snitch_regfile.mem\[418\] i_snitch.i_snitch_regfile.mem\[450\] i_snitch.i_snitch_regfile.mem\[482\]
+ net2974 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_70_790 VPWR VGND sg13g2_fill_2
XFILLER_30_610 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2629 net2851 net3078
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[296\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2643 net2780 net2318 net1318 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[191\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xhold828 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\] VPWR
+ VGND net860 sg13g2_dlygate4sd3_1
Xhold817 i_snitch.i_snitch_regfile.mem\[104\] VPWR VGND net849 sg13g2_dlygate4sd3_1
XFILLER_7_894 VPWR VGND sg13g2_fill_1
XFILLER_6_360 VPWR VGND sg13g2_fill_1
Xhold806 i_snitch.i_snitch_regfile.mem\[473\] VPWR VGND net838 sg13g2_dlygate4sd3_1
Xhold839 i_snitch.i_snitch_regfile.mem\[148\] VPWR VGND net871 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2419 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2585 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xdata_pdata\[14\]_sg13g2_mux2_1_A1 rsp_data_q\[14\] net1035 net3050 data_pdata\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xfanout3270 net3271 net3270 VPWR VGND sg13g2_buf_8
Xfanout3281 net3282 net3281 VPWR VGND sg13g2_buf_8
Xfanout3292 net3300 net3292 VPWR VGND sg13g2_buf_8
Xfanout2580 net2583 net2580 VPWR VGND sg13g2_buf_2
XFILLER_97_687 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[297\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[297\]
+ net3008 i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_a21oi_1_A1_Y net2982 sg13g2_a21oi_1
Xfanout2591 net2592 net2591 VPWR VGND sg13g2_buf_2
XFILLER_69_389 VPWR VGND sg13g2_fill_2
XFILLER_93_860 VPWR VGND sg13g2_decap_8
XFILLER_37_242 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2592 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ net2523 i_snitch.inst_addr_o\[27\] sg13g2_or2_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_80_521 VPWR VGND sg13g2_decap_8
XFILLER_25_426 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q net3278 VGND VPWR i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[326\] clknet_leaf_77_clk sg13g2_dfrbpq_1
XFILLER_80_587 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2448 net2271 net2409 net1165 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[506\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[477\] net2950 VPWR VGND sg13g2_nand2_1
XFILLER_106_203 VPWR VGND sg13g2_decap_8
XFILLER_106_7 VPWR VGND sg13g2_decap_8
XFILLER_88_610 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[14\]_sg13g2_a22oi_1_A1 shift_reg_q\[14\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[14\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A_Y net2827 i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_103_921 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_102_431 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y
+ net2611 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
XFILLER_88_665 VPWR VGND sg13g2_decap_8
XFILLER_57_35 VPWR VGND sg13g2_fill_2
XFILLER_0_569 VPWR VGND sg13g2_decap_8
XFILLER_103_998 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ net1158 VGND sg13g2_inv_1
XFILLER_44_713 VPWR VGND sg13g2_fill_2
XFILLER_28_297 VPWR VGND sg13g2_fill_2
XFILLER_43_256 VPWR VGND sg13g2_decap_8
XFILLER_40_930 VPWR VGND sg13g2_fill_2
XFILLER_11_120 VPWR VGND sg13g2_fill_1
XFILLER_12_632 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_7_135 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B
+ VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B
+ sg13g2_o21ai_1
XFILLER_98_42 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_100_clk clknet_5_18__leaf_clk clknet_leaf_100_clk VPWR VGND sg13g2_buf_8
XFILLER_98_429 VPWR VGND sg13g2_decap_8
XFILLER_105_280 VPWR VGND sg13g2_decap_8
XFILLER_3_385 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2_sg13g2_nor2b_1_Y
+ net3073 net3148 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ VPWR VGND sg13g2_nor2b_2
XFILLER_79_676 VPWR VGND sg13g2_decap_4
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B
+ sg13g2_a21oi_1
XFILLER_93_112 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_66_304 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[346\] clknet_leaf_115_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VGND sg13g2_inv_1
XFILLER_82_808 VPWR VGND sg13g2_fill_2
XFILLER_66_337 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net938 net2445 net2284 VPWR VGND sg13g2_a22oi_1
XFILLER_19_220 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1104 net822 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_75_871 VPWR VGND sg13g2_fill_2
XFILLER_19_242 VPWR VGND sg13g2_fill_1
XFILLER_16_971 VPWR VGND sg13g2_decap_4
XFILLER_35_768 VPWR VGND sg13g2_fill_2
XFILLER_90_896 VPWR VGND sg13g2_decap_8
XFILLER_72_1012 VPWR VGND sg13g2_decap_8
XFILLER_50_727 VPWR VGND sg13g2_fill_2
XFILLER_43_790 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_mux2_1_A1
+ net954 net605 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B
+ i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1 VPWR VGND sg13g2_nand3_1
Xrsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net950 net3063 rsp_data_q\[12\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold603 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\] VPWR
+ VGND net635 sg13g2_dlygate4sd3_1
Xhold614 i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net646 sg13g2_dlygate4sd3_1
Xhold636 i_snitch.sb_q\[2\] VPWR VGND net668 sg13g2_dlygate4sd3_1
Xhold625 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_inv_1_A_Y VPWR VGND net657 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[25\] net1061 net2916 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A_Y net2841 i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xhold647 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\] VPWR
+ VGND net679 sg13g2_dlygate4sd3_1
Xhold669 i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_inv_1_A_Y VPWR VGND net701 sg13g2_dlygate4sd3_1
Xhold658 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_inv_1_A_Y VPWR VGND net690 sg13g2_dlygate4sd3_1
XFILLER_103_217 VPWR VGND sg13g2_decap_8
XFILLER_98_941 VPWR VGND sg13g2_decap_8
Xdata_pdata\[0\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net685 data_pdata\[0\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_100_924 VPWR VGND sg13g2_decap_8
XFILLER_85_613 VPWR VGND sg13g2_fill_2
Xhold1314 i_snitch.inst_addr_o\[24\] VPWR VGND net1346 sg13g2_dlygate4sd3_1
Xhold1325 i_snitch.i_snitch_regfile.mem\[226\] VPWR VGND net1357 sg13g2_dlygate4sd3_1
Xhold1303 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\] VPWR
+ VGND net1335 sg13g2_dlygate4sd3_1
Xhold1358 i_snitch.inst_addr_o\[30\] VPWR VGND net1390 sg13g2_dlygate4sd3_1
Xhold1336 i_snitch.i_snitch_regfile.mem\[229\] VPWR VGND net1368 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[385\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold1347 i_snitch.i_snitch_regfile.mem\[36\] VPWR VGND net1379 sg13g2_dlygate4sd3_1
Xhold1369 i_snitch.inst_addr_o\[28\] VPWR VGND net1401 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2570 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B
+ sg13g2_a21oi_1
XFILLER_80_351 VPWR VGND sg13g2_fill_2
XFILLER_14_919 VPWR VGND sg13g2_fill_2
XFILLER_80_362 VPWR VGND sg13g2_fill_2
XFILLER_41_727 VPWR VGND sg13g2_decap_4
XFILLER_22_952 VPWR VGND sg13g2_decap_8
XFILLER_22_963 VPWR VGND sg13g2_fill_1
XFILLER_40_237 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[273\] VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_nand2_1_B
+ i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_B1 net3164 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_4_105 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[366\] clknet_leaf_85_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net887 net2445 net2252 VPWR VGND sg13g2_a22oi_1
XFILLER_89_930 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D_sg13g2_xor2_1_X
+ net3141 net3144 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D
+ VPWR VGND sg13g2_xor2_1
XFILLER_103_762 VPWR VGND sg13g2_fill_1
XFILLER_103_751 VPWR VGND sg13g2_fill_2
XFILLER_88_440 VPWR VGND sg13g2_fill_1
XFILLER_0_344 VPWR VGND sg13g2_decap_8
XFILLER_1_867 VPWR VGND sg13g2_decap_8
XFILLER_103_795 VPWR VGND sg13g2_decap_8
XFILLER_76_613 VPWR VGND sg13g2_fill_2
XFILLER_102_294 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ net45 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_95_1001 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_A1
+ net1075 VGND sg13g2_inv_1
XFILLER_17_702 VPWR VGND sg13g2_fill_1
XFILLER_90_126 VPWR VGND sg13g2_decap_4
XFILLER_84_690 VPWR VGND sg13g2_decap_8
XFILLER_90_159 VPWR VGND sg13g2_fill_2
XFILLER_56_1018 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_A2
+ VGND VPWR net2569 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C
+ sg13g2_a21oi_1
XFILLER_31_215 VPWR VGND sg13g2_decap_4
XFILLER_32_727 VPWR VGND sg13g2_fill_2
Xi_snitch.inst_addr_o\[26\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[26\]
+ i_snitch.inst_addr_o\[26\] clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_9_978 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_69_7 VPWR VGND sg13g2_fill_1
XFILLER_8_466 VPWR VGND sg13g2_fill_2
XFILLER_4_661 VPWR VGND sg13g2_decap_8
XFILLER_95_966 VPWR VGND sg13g2_decap_8
Xdata_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1 net2683 VPWR data_pdata\[31\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[31\]_sg13g2_a21oi_1_A2_Y net3069 sg13g2_o21ai_1
XFILLER_63_852 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[112\]
+ net2997 i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_req_register.data_o\[45\]_sg13g2_o21ai_1_Y i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.data_o\[45\] VGND net3169 i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_23_749 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[386\] clknet_leaf_13_clk sg13g2_dfrbpq_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_95_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[175\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[175\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net906 net2678 net2775 VPWR VGND sg13g2_a22oi_1
Xhold400 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\] VPWR
+ VGND net432 sg13g2_dlygate4sd3_1
Xhold411 strb_reg_q\[5\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold433 shift_reg_q\[4\] VPWR VGND net465 sg13g2_dlygate4sd3_1
Xhold422 i_snitch.i_snitch_regfile.mem\[446\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold444 shift_reg_q\[13\] VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold477 shift_reg_q\[18\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold455 shift_reg_q\[14\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold466 shift_reg_q\[19\] VPWR VGND net498 sg13g2_dlygate4sd3_1
XFILLER_1_119 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2557 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xhold499 i_snitch.sb_q\[8\] VPWR VGND net531 sg13g2_dlygate4sd3_1
Xhold488 shift_reg_q\[11\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net520 sg13g2_dlygate4sd3_1
Xhold1100 i_snitch.i_snitch_regfile.mem\[213\] VPWR VGND net1132 sg13g2_dlygate4sd3_1
XFILLER_86_944 VPWR VGND sg13g2_decap_8
Xhold1122 rsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1154
+ sg13g2_dlygate4sd3_1
Xhold1111 i_snitch.i_snitch_regfile.mem\[275\] VPWR VGND net1143 sg13g2_dlygate4sd3_1
Xhold1133 i_snitch.i_snitch_regfile.mem\[115\] VPWR VGND net1165 sg13g2_dlygate4sd3_1
XFILLER_100_765 VPWR VGND sg13g2_fill_1
XFILLER_85_476 VPWR VGND sg13g2_fill_1
XFILLER_79_1007 VPWR VGND sg13g2_decap_8
Xhold1155 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] VPWR
+ VGND net1187 sg13g2_dlygate4sd3_1
Xhold1144 i_snitch.i_snitch_regfile.mem\[411\] VPWR VGND net1176 sg13g2_dlygate4sd3_1
Xhold1166 i_snitch.i_snitch_regfile.mem\[48\] VPWR VGND net1198 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[484\]_sg13g2_nor3_1_A net1313 net2855 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_100_798 VPWR VGND sg13g2_decap_8
XFILLER_85_498 VPWR VGND sg13g2_fill_1
Xhold1188 i_snitch.i_snitch_regfile.mem\[405\] VPWR VGND net1220 sg13g2_dlygate4sd3_1
Xhold1199 i_snitch.i_snitch_regfile.mem\[302\] VPWR VGND net1231 sg13g2_dlygate4sd3_1
Xhold1177 i_snitch.i_snitch_regfile.mem\[294\] VPWR VGND net1209 sg13g2_dlygate4sd3_1
XFILLER_38_370 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y net2723
+ net3148 VPWR VGND sg13g2_a22oi_1
XFILLER_14_705 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[205\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_54_58 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2590 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A
+ sg13g2_or2_1
XFILLER_9_208 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_103_1005 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1
+ net770 net569 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2414
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_436 VPWR VGND sg13g2_decap_8
XFILLER_10_999 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_nor3_1_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ net76 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ VPWR VGND sg13g2_nor3_2
XFILLER_1_664 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_88_281 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_nand2b_1_A_N_Y
+ net3027 i_snitch.i_snitch_regfile.mem\[91\] VPWR VGND sg13g2_nand2b_1
XFILLER_77_977 VPWR VGND sg13g2_decap_8
XFILLER_49_668 VPWR VGND sg13g2_fill_2
XFILLER_48_167 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2831
+ VPWR i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_1_Y
+ sg13g2_o21ai_1
Xshift_reg_q\[7\]_sg13g2_nor2_1_A net492 net2731 shift_reg_q\[7\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_92_969 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[501\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[501\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2268 net2367 net1189 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[125\]
+ net2998 i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_1 i_snitch.i_snitch_regfile.mem\[120\]
+ net2807 i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_1_Y VPWR VGND sg13g2_nor2_1
XFILLER_45_841 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2866
+ net2660 VPWR VGND sg13g2_nand2_1
XFILLER_72_660 VPWR VGND sg13g2_fill_1
XFILLER_17_587 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2361 net1079 net2680 net2769 VPWR VGND sg13g2_a22oi_1
XFILLER_9_720 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1365 net3065 rsp_data_q\[1\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xor2_1
XFILLER_67_4 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[502\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[502\]
+ net3135 i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
XFILLER_8_274 VPWR VGND sg13g2_decap_4
XFILLER_5_970 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_101_529 VPWR VGND sg13g2_fill_1
XFILLER_101_518 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[225\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_95_752 VPWR VGND sg13g2_decap_8
XFILLER_95_730 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_q\[2\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[2\] i_snitch.sb_q\[2\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_83_914 VPWR VGND sg13g2_decap_8
XFILLER_94_295 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ net103 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1297 net2495 net1187 VPWR VGND sg13g2_a22oi_1
XFILLER_27_329 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N
+ net2751 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_63_682 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B
+ net2631 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2639 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_10_218 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2457 net2855 i_snitch.i_snitch_regfile.mem\[484\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
XFILLER_85_1011 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[255\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2328
+ sg13g2_o21ai_1
XFILLER_104_301 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2885
+ net2661 VPWR VGND sg13g2_nand2_1
XFILLER_105_868 VPWR VGND sg13g2_decap_8
Xfanout2409 net2410 net2409 VPWR VGND sg13g2_buf_8
XFILLER_104_378 VPWR VGND sg13g2_decap_8
XFILLER_105_42 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2 VPWR VGND i_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_B2
+ i_snitch.pc_d\[12\]_sg13g2_mux2_1_A1_X i_snitch.pc_d\[22\] i_snitch.pc_d\[16\] i_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1 sg13g2_a221oi_1
XFILLER_74_903 VPWR VGND sg13g2_fill_1
XFILLER_59_999 VPWR VGND sg13g2_fill_2
XFILLER_85_273 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_mux2_1_A0_X net3103 net2826 i_snitch.i_snitch_regfile.mem\[63\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2360 net812 net2646 net2767 VPWR VGND sg13g2_a22oi_1
XFILLER_46_627 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2535 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_A sg13g2_a21oi_1
XFILLER_65_68 VPWR VGND sg13g2_fill_1
XFILLER_26_340 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_92_1004 VPWR VGND sg13g2_decap_8
XFILLER_14_513 VPWR VGND sg13g2_fill_1
XFILLER_60_129 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_80_clk clknet_5_28__leaf_clk clknet_leaf_80_clk VPWR VGND sg13g2_buf_8
XFILLER_26_395 VPWR VGND sg13g2_decap_4
XFILLER_41_310 VPWR VGND sg13g2_fill_2
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[245\] clknet_leaf_98_clk sg13g2_dfrbpq_1
Xrebuffer382 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y
+ net414 VPWR VGND sg13g2_buf_1
XFILLER_5_244 VPWR VGND sg13g2_fill_1
Xfanout2921 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_A2 net2921 VPWR
+ VGND sg13g2_buf_8
Xfanout2910 data_pdata\[19\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2910 VPWR VGND
+ sg13g2_buf_8
Xfanout2932 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net2932 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3042
+ net2649 VPWR VGND sg13g2_nand2_1
Xfanout2954 net2955 net2954 VPWR VGND sg13g2_buf_8
Xfanout2943 net2945 net2943 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C
+ net2848 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_77_730 VPWR VGND sg13g2_fill_1
Xfanout2965 net2966 net2965 VPWR VGND sg13g2_buf_8
Xfanout2998 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2998 VPWR VGND sg13g2_buf_8
XFILLER_7_1011 VPWR VGND sg13g2_decap_8
Xfanout2987 net2989 net2987 VPWR VGND sg13g2_buf_8
Xfanout2976 net2996 net2976 VPWR VGND sg13g2_buf_8
Xrsp_data_q\[9\]_sg13g2_dfrbpq_1_Q net3239 VGND VPWR rsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[9\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] net582 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_37_649 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1381 net2493 net1213 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ VGND net2572 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_92_755 VPWR VGND sg13g2_decap_8
XFILLER_80_917 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_C
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B_X
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2_Y VPWR VGND sg13g2_and3_1
XFILLER_65_969 VPWR VGND sg13g2_decap_4
XFILLER_18_852 VPWR VGND sg13g2_fill_2
XFILLER_52_619 VPWR VGND sg13g2_decap_4
XFILLER_51_118 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3094 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
Xclkbuf_leaf_71_clk clknet_5_24__leaf_clk clknet_leaf_71_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2357
+ sg13g2_o21ai_1
XFILLER_20_527 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.inst_addr_o\[25\] net2523 VPWR VGND sg13g2_xnor2_1
XFILLER_9_583 VPWR VGND sg13g2_fill_2
XFILLER_9_572 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[45\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X
+ net2510 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net929 net2451 net2271 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
XFILLER_99_365 VPWR VGND sg13g2_decap_8
XFILLER_102_849 VPWR VGND sg13g2_decap_8
XFILLER_101_315 VPWR VGND sg13g2_decap_8
XFILLER_59_229 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_19_17 VPWR VGND sg13g2_fill_1
XFILLER_68_774 VPWR VGND sg13g2_fill_2
XFILLER_68_763 VPWR VGND sg13g2_decap_8
XFILLER_83_744 VPWR VGND sg13g2_decap_8
XFILLER_55_446 VPWR VGND sg13g2_decap_8
XFILLER_83_788 VPWR VGND sg13g2_fill_1
XFILLER_70_449 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_62_clk clknet_5_29__leaf_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q net3251 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[9\] clknet_leaf_18_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[265\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_24_844 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_24_888 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q
+ net3238 VGND VPWR net1004 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net3134 net2851 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1
+ net2629 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2862
+ net2653 VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1297 net3066 rsp_data_q\[10\] VPWR VGND sg13g2_a22oi_1
XFILLER_13_1027 VPWR VGND sg13g2_fill_2
XFILLER_100_1008 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[356\]_sg13g2_nor3_1_A net1284 net2879 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[356\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_2_203 VPWR VGND sg13g2_fill_1
Xfanout2239 net2239 net68 VPWR VGND sg13g2_buf_16
XFILLER_104_175 VPWR VGND sg13g2_decap_8
XFILLER_78_538 VPWR VGND sg13g2_fill_1
XFILLER_59_730 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2578 sg13g2_a21oi_1
XFILLER_101_882 VPWR VGND sg13g2_decap_8
XFILLER_86_571 VPWR VGND sg13g2_fill_1
XFILLER_59_796 VPWR VGND sg13g2_decap_8
XFILLER_47_925 VPWR VGND sg13g2_fill_1
XFILLER_19_616 VPWR VGND sg13g2_fill_2
XFILLER_18_126 VPWR VGND sg13g2_fill_2
XFILLER_61_405 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2539 sg13g2_a21oi_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y
+ net3078 net2537 i_snitch.inst_addr_o\[10\] i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_53_clk clknet_5_26__leaf_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
XFILLER_14_365 VPWR VGND sg13g2_decap_8
XFILLER_14_376 VPWR VGND sg13g2_fill_2
XFILLER_30_825 VPWR VGND sg13g2_decap_8
XFILLER_42_685 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_69_505 VPWR VGND sg13g2_fill_1
Xfanout2751 net2754 net2751 VPWR VGND sg13g2_buf_8
Xfanout2762 net2763 net2762 VPWR VGND sg13g2_buf_2
Xfanout2740 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2740 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2742
+ net2656 VPWR VGND sg13g2_nand2_1
XFILLER_2_53 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[285\] clknet_leaf_95_clk sg13g2_dfrbpq_1
Xfanout2784 net2785 net2784 VPWR VGND sg13g2_buf_8
Xfanout2795 net2799 net2795 VPWR VGND sg13g2_buf_8
Xfanout2773 net2776 net2773 VPWR VGND sg13g2_buf_8
XFILLER_77_571 VPWR VGND sg13g2_fill_1
XFILLER_92_552 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR net776 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q
+ net3185 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
XFILLER_92_585 VPWR VGND sg13g2_fill_1
XFILLER_80_769 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_44_clk clknet_5_15__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_60_482 VPWR VGND sg13g2_fill_2
XFILLER_21_836 VPWR VGND sg13g2_fill_1
Xdata_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[12\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[28\]_sg13g2_nand2b_1_B_Y net3152 data_pdata\[20\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[12\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
XFILLER_21_858 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A
+ net3080 net2851 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2481 net2421 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y
+ net2500 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[209\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[209\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2339 net1039 net2664 net2793 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nand2b_1_A_N_Y
+ net3026 i_snitch.i_snitch_regfile.mem\[69\] VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2786
+ net2694 VPWR VGND sg13g2_nand2_1
XFILLER_99_140 VPWR VGND sg13g2_decap_8
XFILLER_82_1014 VPWR VGND sg13g2_decap_8
XFILLER_101_112 VPWR VGND sg13g2_decap_8
XFILLER_88_847 VPWR VGND sg13g2_decap_8
XFILLER_87_335 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2
+ net2955 net2752 net3089 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[104\] clknet_leaf_71_clk sg13g2_dfrbpq_1
XFILLER_102_679 VPWR VGND sg13g2_fill_2
XFILLER_102_668 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B_sg13g2_nor2_1_Y
+ net3085 net3087 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B
+ VPWR VGND sg13g2_nor2_2
XFILLER_101_189 VPWR VGND sg13g2_decap_8
XFILLER_96_880 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2544 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ net2612 VPWR VGND sg13g2_a22oi_1
XFILLER_102_21 VPWR VGND sg13g2_decap_8
XFILLER_71_725 VPWR VGND sg13g2_fill_2
XFILLER_71_714 VPWR VGND sg13g2_decap_4
XFILLER_16_619 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_15_129 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_35_clk clknet_5_8__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_71_769 VPWR VGND sg13g2_fill_1
XFILLER_52_972 VPWR VGND sg13g2_fill_2
XFILLER_24_663 VPWR VGND sg13g2_fill_1
XFILLER_102_98 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2720 i_snitch.inst_addr_o\[29\] sg13g2_a21oi_2
XFILLER_11_357 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0 net3137 i_snitch.i_snitch_regfile.mem\[152\]
+ i_snitch.i_snitch_regfile.mem\[184\] i_snitch.i_snitch_regfile.mem\[216\] i_snitch.i_snitch_regfile.mem\[248\]
+ net3111 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_106_941 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B
+ net2579 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2467 net2262 net2389 net1225 VPWR VGND sg13g2_a22oi_1
XFILLER_79_869 VPWR VGND sg13g2_decap_4
XFILLER_4_1025 VPWR VGND sg13g2_decap_4
Xdata_pdata\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C net3149 data_pdata\[13\]_sg13g2_nor2b_1_A_Y
+ data_pdata\[5\]_sg13g2_nor2_1_B_Y data_pdata\[5\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_19_435 VPWR VGND sg13g2_fill_1
XFILLER_74_563 VPWR VGND sg13g2_fill_1
XFILLER_46_287 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_26_clk clknet_5_8__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_99_7 VPWR VGND sg13g2_decap_8
XFILLER_43_983 VPWR VGND sg13g2_fill_1
XFILLER_14_162 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[264\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_B1
+ net990 net2306 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[124\] clknet_leaf_99_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2449
+ net2514 net2902 net2868 VPWR VGND sg13g2_a22oi_1
Xhold807 i_snitch.i_snitch_regfile.mem\[364\] VPWR VGND net839 sg13g2_dlygate4sd3_1
XFILLER_10_390 VPWR VGND sg13g2_fill_2
Xhold818 i_snitch.i_snitch_regfile.mem\[397\] VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold829 i_snitch.i_snitch_regfile.mem\[32\] VPWR VGND net861 sg13g2_dlygate4sd3_1
XFILLER_97_600 VPWR VGND sg13g2_fill_2
Xfanout3260 net3261 net3260 VPWR VGND sg13g2_buf_8
Xi_req_arb.data_i\[43\]_sg13g2_dfrbpq_1_Q net3305 VGND VPWR i_snitch.pc_d\[8\] i_req_arb.data_i\[43\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_2
Xfanout3271 net3272 net3271 VPWR VGND sg13g2_buf_8
Xfanout3282 net3329 net3282 VPWR VGND sg13g2_buf_8
Xfanout2581 net2583 net2581 VPWR VGND sg13g2_buf_8
XFILLER_97_666 VPWR VGND sg13g2_decap_8
Xfanout2570 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X
+ net2570 VPWR VGND sg13g2_buf_8
XFILLER_85_806 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[23\]_sg13g2_dfrbpq_1_Q net3199 VGND VPWR net512 shift_reg_q\[23\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
Xfanout3293 net3294 net3293 VPWR VGND sg13g2_buf_8
Xfanout2592 net2593 net2592 VPWR VGND sg13g2_buf_8
XFILLER_57_519 VPWR VGND sg13g2_decap_4
XFILLER_38_722 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_37_210 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[91\]
+ i_snitch.i_snitch_regfile.mem\[123\] net3119 i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_38_788 VPWR VGND sg13g2_fill_2
XFILLER_92_382 VPWR VGND sg13g2_fill_2
XFILLER_65_596 VPWR VGND sg13g2_decap_8
XFILLER_19_980 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_17_clk clknet_5_13__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_18_490 VPWR VGND sg13g2_decap_8
XFILLER_21_622 VPWR VGND sg13g2_fill_1
XFILLER_21_655 VPWR VGND sg13g2_fill_1
XFILLER_33_493 VPWR VGND sg13g2_fill_1
XFILLER_21_666 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1 i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_X net3096 i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VPWR VGND
+ sg13g2_a22oi_1
XFILLER_20_176 VPWR VGND sg13g2_fill_2
Xrsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1381 net3066 net8 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0 net124 i_snitch.i_snitch_regfile.mem\[390\]
+ i_snitch.i_snitch_regfile.mem\[422\] i_snitch.i_snitch_regfile.mem\[454\] i_snitch.i_snitch_regfile.mem\[486\]
+ net3107 i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_106_259 VPWR VGND sg13g2_decap_8
XFILLER_103_900 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C i_snitch.inst_addr_o\[31\]
+ net2303 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_103_977 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B
+ net2959 i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_88_699 VPWR VGND sg13g2_decap_8
XFILLER_87_176 VPWR VGND sg13g2_fill_2
XFILLER_87_165 VPWR VGND sg13g2_fill_1
XFILLER_57_58 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[412\] VGND sg13g2_inv_1
XFILLER_75_338 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[249\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[249\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net1006 net2438 net2266 VPWR VGND sg13g2_a22oi_1
XFILLER_56_574 VPWR VGND sg13g2_fill_2
XFILLER_44_703 VPWR VGND sg13g2_fill_1
XFILLER_73_46 VPWR VGND sg13g2_decap_4
XFILLER_56_596 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[144\] clknet_leaf_90_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[228\]_sg13g2_nor3_1_A net1338 net2874 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_32_909 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_43_279 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_419 VPWR VGND sg13g2_decap_8
XFILLER_106_1025 VPWR VGND sg13g2_decap_4
XFILLER_52_791 VPWR VGND sg13g2_decap_4
XFILLER_11_143 VPWR VGND sg13g2_decap_8
XFILLER_8_659 VPWR VGND sg13g2_decap_8
XFILLER_99_909 VPWR VGND sg13g2_decap_8
XFILLER_98_21 VPWR VGND sg13g2_decap_8
Xdata_pdata\[30\]_sg13g2_a21oi_1_A2 VGND VPWR net3162 data_pdata\[30\] data_pdata\[30\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[22\]_sg13g2_nor2b_1_B_N_Y sg13g2_a21oi_1
XFILLER_98_98 VPWR VGND sg13g2_decap_8
XFILLER_79_633 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[446\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_26_1026 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[481\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net447 net2368 VPWR VGND sg13g2_nand2_1
XFILLER_67_839 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y
+ net2762 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 net2852 net3090
+ VPWR VGND sg13g2_a22oi_1
XFILLER_93_179 VPWR VGND sg13g2_fill_1
XFILLER_81_319 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[440\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2383 net796 net2665 net2863 VPWR VGND sg13g2_a22oi_1
XFILLER_47_596 VPWR VGND sg13g2_fill_2
XFILLER_34_202 VPWR VGND sg13g2_decap_8
XFILLER_90_875 VPWR VGND sg13g2_decap_8
XFILLER_16_950 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net3038 net2905 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2697 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_Y VPWR VGND sg13g2_nand2_1
XFILLER_72_1002 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net907 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] net2913
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_452 VPWR VGND sg13g2_decap_8
XFILLER_8_63 VPWR VGND sg13g2_fill_2
Xhold604 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net636 sg13g2_dlygate4sd3_1
Xhold626 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\] VPWR
+ VGND net658 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_a22oi_1_B2_Y
+ net2324 net704 net2689 net2895 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B
+ net2499 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xhold615 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\] VPWR
+ VGND net647 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1
+ net2637 i_req_arb.data_i\[43\] i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ net2722 sg13g2_a221oi_1
Xhold637 i_snitch.inst_addr_o\[1\] VPWR VGND net669 sg13g2_dlygate4sd3_1
Xhold659 i_snitch.i_snitch_regfile.mem\[277\] VPWR VGND net691 sg13g2_dlygate4sd3_1
Xhold648 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net680 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_5_2__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_98_920 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0 net3124 i_snitch.i_snitch_regfile.mem\[159\]
+ i_snitch.i_snitch_regfile.mem\[191\] i_snitch.i_snitch_regfile.mem\[223\] i_snitch.i_snitch_regfile.mem\[255\]
+ net3103 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
XFILLER_100_903 VPWR VGND sg13g2_decap_8
Xfanout3090 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_X
+ net3090 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[164\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[164\] clknet_leaf_13_clk sg13g2_dfrbpq_1
XFILLER_98_997 VPWR VGND sg13g2_decap_8
Xhold1304 rsp_data_q\[10\] VPWR VGND net1336 sg13g2_dlygate4sd3_1
Xhold1315 rsp_data_q\[25\] VPWR VGND net1347 sg13g2_dlygate4sd3_1
XFILLER_58_828 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2606 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_97_496 VPWR VGND sg13g2_fill_2
Xhold1337 rsp_data_q\[2\] VPWR VGND net1369 sg13g2_dlygate4sd3_1
XFILLER_69_198 VPWR VGND sg13g2_fill_2
Xhold1359 i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q VPWR VGND
+ net1391 sg13g2_dlygate4sd3_1
Xhold1348 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\] VPWR
+ VGND net1380 sg13g2_dlygate4sd3_1
Xhold1326 i_snitch.i_snitch_regfile.mem\[98\] VPWR VGND net1358 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y
+ i_snitch.sb_q\[3\] net2803 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_27_39 VPWR VGND sg13g2_fill_1
XFILLER_25_213 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_81_886 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A
+ VPWR i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A_Y
+ net441 VGND sg13g2_inv_1
XFILLER_53_577 VPWR VGND sg13g2_fill_2
XFILLER_40_216 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[460\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[460\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net762 net2691 net2741 VPWR VGND sg13g2_a22oi_1
Xi_req_register.data_o\[5\]_sg13g2_inv_1_A_Y_sg13g2_nor2_1_B net3053 i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y
+ cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 VPWR VGND sg13g2_nor2_2
XFILLER_88_430 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0 net3133 i_snitch.i_snitch_regfile.mem\[278\]
+ i_snitch.i_snitch_regfile.mem\[310\] i_snitch.i_snitch_regfile.mem\[342\] i_snitch.i_snitch_regfile.mem\[374\]
+ net3113 i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_1_846 VPWR VGND sg13g2_decap_8
XFILLER_103_774 VPWR VGND sg13g2_decap_8
XFILLER_89_986 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_fill_2
XFILLER_102_273 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_84_34 VPWR VGND sg13g2_decap_8
XFILLER_29_552 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B
+ net2590 sg13g2_or2_1
XFILLER_91_639 VPWR VGND sg13g2_decap_4
XFILLER_1_1028 VPWR VGND sg13g2_fill_1
XFILLER_29_596 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y i_snitch.pc_d\[11\] i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2 net2307 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_71_341 VPWR VGND sg13g2_decap_4
Xdata_pdata\[17\]_sg13g2_nor2b_1_B_N net3156 data_pdata\[17\] data_pdata\[17\]_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_Y
+ VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ VGND net46 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y
+ sg13g2_o21ai_1
XFILLER_13_931 VPWR VGND sg13g2_fill_1
XFILLER_13_953 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[289\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2901 net2779 net2317 net1316 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_A
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nor4_1
Xrsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1306 net3065 net1183 VPWR VGND sg13g2_a22oi_1
XFILLER_9_968 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[184\] clknet_leaf_57_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1
+ net2705 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_79_430 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0 net3130 i_snitch.i_snitch_regfile.mem\[397\]
+ i_snitch.i_snitch_regfile.mem\[429\] i_snitch.i_snitch_regfile.mem\[461\] i_snitch.i_snitch_regfile.mem\[493\]
+ net3109 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q net3257 VGND VPWR i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[32\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_95_945 VPWR VGND sg13g2_decap_8
Xdata_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2681 data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_81_116 VPWR VGND sg13g2_fill_1
XFILLER_63_820 VPWR VGND sg13g2_decap_8
XFILLER_48_883 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y net3004 sg13g2_o21ai_1
XFILLER_35_500 VPWR VGND sg13g2_fill_1
XFILLER_62_341 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[319\] clknet_leaf_70_clk sg13g2_dfrbpq_1
XFILLER_23_706 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2410 net1015 net2692 net2869 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_nor3_1_A net1289 net2886 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nor2b_1
XFILLER_50_558 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[2\]_sg13g2_dfrbpq_1_Q net3185 VGND VPWR net518 strb_reg_q\[2\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
XFILLER_88_0 VPWR VGND sg13g2_fill_2
Xstrb_reg_q\[5\]_sg13g2_nor2_1_A strb_reg_q\[5\] net2727 strb_reg_q\[5\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xdata_pdata\[25\]_sg13g2_mux2_1_A1 rsp_data_q\[25\] net945 net3048 data_pdata\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net3144 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[480\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2367 net973 net2903 net2855 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[30\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[30\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[30\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_and2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net3082 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ net2850 net3074 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ net2754 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2377
+ sg13g2_o21ai_1
Xhold401 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net433 sg13g2_dlygate4sd3_1
XFILLER_8_990 VPWR VGND sg13g2_decap_8
Xhold434 shift_reg_q\[4\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net466 sg13g2_dlygate4sd3_1
Xhold445 shift_reg_q\[13\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold423 i_snitch.i_snitch_regfile.mem\[430\] VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold412 i_snitch.i_snitch_regfile.mem\[225\] VPWR VGND net444 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q
+ net3231 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xhold467 shift_reg_q\[19\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold456 i_snitch.sb_q\[4\] VPWR VGND net488 sg13g2_dlygate4sd3_1
Xhold478 i_snitch.i_snitch_regfile.mem\[442\] VPWR VGND net510 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold489 shift_reg_q\[3\] VPWR VGND net521 sg13g2_dlygate4sd3_1
XFILLER_86_923 VPWR VGND sg13g2_decap_8
XFILLER_85_411 VPWR VGND sg13g2_decap_8
XFILLER_58_603 VPWR VGND sg13g2_decap_4
XFILLER_57_102 VPWR VGND sg13g2_fill_1
Xhold1101 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] VPWR
+ VGND net1133 sg13g2_dlygate4sd3_1
XFILLER_58_647 VPWR VGND sg13g2_decap_8
Xhold1123 i_snitch.i_snitch_regfile.mem\[414\] VPWR VGND net1155 sg13g2_dlygate4sd3_1
Xhold1112 i_snitch.i_snitch_regfile.mem\[237\] VPWR VGND net1144 sg13g2_dlygate4sd3_1
XFILLER_73_617 VPWR VGND sg13g2_fill_1
Xhold1134 i_snitch.inst_addr_o\[19\] VPWR VGND net1166 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2385
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand2_2
Xhold1145 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\] VPWR
+ VGND net1177 sg13g2_dlygate4sd3_1
Xhold1156 i_snitch.i_snitch_regfile.mem\[185\] VPWR VGND net1188 sg13g2_dlygate4sd3_1
Xhold1167 i_snitch.i_snitch_regfile.mem\[505\] VPWR VGND net1199 sg13g2_dlygate4sd3_1
XFILLER_54_831 VPWR VGND sg13g2_fill_1
Xhold1189 i_snitch.i_snitch_regfile.mem\[309\] VPWR VGND net1221 sg13g2_dlygate4sd3_1
Xhold1178 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] VPWR
+ VGND net1210 sg13g2_dlygate4sd3_1
XFILLER_54_37 VPWR VGND sg13g2_decap_4
XFILLER_53_374 VPWR VGND sg13g2_fill_1
XFILLER_41_514 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[510\] clknet_leaf_93_clk sg13g2_dfrbpq_1
XFILLER_13_249 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_41_547 VPWR VGND sg13g2_fill_1
XFILLER_41_558 VPWR VGND sg13g2_fill_1
Xdata_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1 net2682 VPWR data_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[25\]_sg13g2_a21oi_1_A2_Y net3069 sg13g2_o21ai_1
XFILLER_103_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y
+ i_snitch.sb_q\[2\] net3122 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_905 VPWR VGND sg13g2_fill_1
XFILLER_10_967 VPWR VGND sg13g2_fill_1
Xdata_pdata\[27\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[27\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[27\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[52\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_6_949 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2735 shift_reg_q\[12\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[8\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[8\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_1_643 VPWR VGND sg13g2_decap_8
Xhold990 i_snitch.i_snitch_regfile.mem\[381\] VPWR VGND net1022 sg13g2_dlygate4sd3_1
XFILLER_103_571 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[13\]_sg13g2_xnor2_1_A i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A
+ i_snitch.inst_addr_o\[13\] net2528 VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[339\] clknet_leaf_116_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net694 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2387 net3038 i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D net2909
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2352 net741 net2903 net2887 VPWR VGND sg13g2_a22oi_1
XFILLER_23_1018 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2596 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_92_948 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_o21ai_1_A1 net3018 VPWR i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[48\] net2987 sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2417 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[269\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_60_878 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[27\]_sg13g2_a22oi_1_A1 shift_reg_q\[27\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[27\] VPWR VGND sg13g2_a22oi_1
XFILLER_81_7 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_2
XFILLER_9_754 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[129\]
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_Y
+ net3013 sg13g2_a21oi_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ net122 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_req_arb.data_i\[39\] sg13g2_a21oi_1
XFILLER_9_787 VPWR VGND sg13g2_decap_8
XFILLER_12_282 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A_X
+ VPWR VGND sg13g2_or3_1
XFILLER_99_503 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand4_1_A
+ net2927 net3036 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_A
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ sg13g2_nand4_1
XFILLER_5_53 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 i_req_arb.data_i\[39\] VPWR
+ VGND sg13g2_nand2b_1
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1
+ i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_95_786 VPWR VGND sg13g2_decap_8
XFILLER_94_252 VPWR VGND sg13g2_fill_2
XFILLER_68_989 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_82_436 VPWR VGND sg13g2_fill_2
XFILLER_82_425 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[72\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_24_18 VPWR VGND sg13g2_fill_2
XFILLER_51_889 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[359\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2450 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_A_N
+ VGND net2750 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net871 net2671 net2888 VPWR VGND sg13g2_a22oi_1
XFILLER_2_418 VPWR VGND sg13g2_fill_1
XFILLER_2_429 VPWR VGND sg13g2_fill_1
XFILLER_105_847 VPWR VGND sg13g2_decap_8
XFILLER_104_357 VPWR VGND sg13g2_decap_8
XFILLER_105_21 VPWR VGND sg13g2_decap_8
XFILLER_100_563 VPWR VGND sg13g2_decap_4
XFILLER_100_541 VPWR VGND sg13g2_decap_4
XFILLER_19_809 VPWR VGND sg13g2_fill_2
XFILLER_105_98 VPWR VGND sg13g2_decap_8
XFILLER_86_797 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y
+ net2524 VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A
+ VGND i_snitch.inst_addr_o\[29\] i_snitch.inst_addr_o\[30\] sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2509 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1
+ net2302 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_27_875 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_42_889 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1
+ net1003 net576 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.inst_addr_o\[19\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.pc_d\[19\]
+ i_snitch.inst_addr_o\[19\] clknet_leaf_53_clk sg13g2_dfrbpq_2
XFILLER_41_377 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ VGND net2704 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ net49 net2515 VPWR VGND sg13g2_nand2_2
Xi_req_register.data_o\[5\]_sg13g2_inv_1_A i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y
+ i_req_register.data_o\[5\] VPWR VGND sg13g2_inv_2
XFILLER_10_797 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3059 net1382 net3064 net6 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1 net2762
+ VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_5_289 VPWR VGND sg13g2_decap_8
Xfanout2911 data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2911 VPWR VGND
+ sg13g2_buf_8
Xfanout2900 data_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2900 VPWR
+ VGND sg13g2_buf_8
Xfanout2922 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D
+ net2922 VPWR VGND sg13g2_buf_8
Xfanout2955 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ net2955 VPWR VGND sg13g2_buf_8
Xfanout2944 net2945 net2944 VPWR VGND sg13g2_buf_8
XFILLER_2_985 VPWR VGND sg13g2_decap_8
Xfanout2933 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2
+ net2933 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ net2585 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ net2591 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xfanout2966 net2967 net2966 VPWR VGND sg13g2_buf_8
XFILLER_49_422 VPWR VGND sg13g2_decap_4
Xfanout2977 net2979 net2977 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[92\] clknet_leaf_101_clk sg13g2_dfrbpq_1
Xfanout2988 net2989 net2988 VPWR VGND sg13g2_buf_8
Xfanout2999 net3003 net2999 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q
+ net3240 VGND VPWR net771 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_B_N
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_92_789 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[379\] clknet_leaf_115_clk sg13g2_dfrbpq_1
XFILLER_44_160 VPWR VGND sg13g2_fill_2
XFILLER_33_845 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[168\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2343 net953 net2643 net2773 VPWR VGND sg13g2_a22oi_1
XFILLER_60_697 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[88\]_sg13g2_o21ai_1_A1 net3111 VPWR i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[88\] net3138 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2639 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_99_311 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y
+ net434 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2363
+ sg13g2_o21ai_1
XFILLER_102_828 VPWR VGND sg13g2_decap_8
XFILLER_87_506 VPWR VGND sg13g2_fill_1
XFILLER_67_252 VPWR VGND sg13g2_fill_2
XFILLER_95_583 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2697 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B
+ net2541 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2393
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_X
+ net3092 net2929 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_27_149 VPWR VGND sg13g2_decap_8
XFILLER_70_417 VPWR VGND sg13g2_decap_4
XFILLER_35_39 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1
+ net2684 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_Y
+ VGND net2848 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2
+ sg13g2_o21ai_1
XFILLER_51_653 VPWR VGND sg13g2_fill_1
XFILLER_23_333 VPWR VGND sg13g2_fill_2
XFILLER_23_388 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2276
+ sg13g2_o21ai_1
XFILLER_105_622 VPWR VGND sg13g2_fill_1
XFILLER_105_688 VPWR VGND sg13g2_fill_1
XFILLER_105_677 VPWR VGND sg13g2_decap_8
XFILLER_104_154 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X net3096 i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VPWR VGND
+ sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[399\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[360\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[360\]
+ net3133 i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2450
+ net2262 net2667 net2870 VPWR VGND sg13g2_a22oi_1
XFILLER_101_861 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2605 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_93_509 VPWR VGND sg13g2_decap_8
XFILLER_59_742 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[188\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[188\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2443 net2246 net2342 net1190 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ net2587 VPWR VGND sg13g2_a22oi_1
XFILLER_74_734 VPWR VGND sg13g2_fill_2
XFILLER_74_767 VPWR VGND sg13g2_fill_1
XFILLER_73_211 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D
+ net764 VGND sg13g2_inv_1
XFILLER_46_447 VPWR VGND sg13g2_decap_8
XFILLER_92_67 VPWR VGND sg13g2_fill_1
Xrebuffer90 net2536 net122 VPWR VGND sg13g2_buf_1
XFILLER_70_973 VPWR VGND sg13g2_fill_1
XFILLER_15_856 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_mux2_1_A0_X net3103 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a22oi_1_A1_A2
+ i_snitch.i_snitch_regfile.mem\[36\] VPWR VGND sg13g2_a22oi_1
XFILLER_41_174 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0
+ VGND net2701 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1
+ net488 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
XFILLER_6_510 VPWR VGND sg13g2_fill_2
XFILLER_10_594 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[96\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_nand2b_1_A_N_Y
+ net2983 i_snitch.i_snitch_regfile.mem\[96\] VPWR VGND sg13g2_nand2b_1
XFILLER_29_1024 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1 VPWR VGND
+ net2933 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y net3089 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[218\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\] VGND sg13g2_inv_1
Xfanout2730 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y net2730
+ VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[37\]
+ net2824 i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1_Y net2821 sg13g2_a21oi_1
XFILLER_97_859 VPWR VGND sg13g2_decap_8
XFILLER_96_314 VPWR VGND sg13g2_decap_8
Xfanout2752 net2754 net2752 VPWR VGND sg13g2_buf_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B
+ net2848 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xfanout2763 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_Y
+ net2763 VPWR VGND sg13g2_buf_8
Xfanout2741 net2743 net2741 VPWR VGND sg13g2_buf_8
XFILLER_2_782 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X net2302 net1196 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[7\] VPWR VGND sg13g2_a21o_1
XFILLER_2_32 VPWR VGND sg13g2_decap_8
Xfanout2774 net2776 net2774 VPWR VGND sg13g2_buf_8
Xfanout2796 net2799 net2796 VPWR VGND sg13g2_buf_8
Xfanout2785 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X
+ net2785 VPWR VGND sg13g2_buf_8
XFILLER_80_726 VPWR VGND sg13g2_fill_1
XFILLER_80_715 VPWR VGND sg13g2_decap_4
XFILLER_65_778 VPWR VGND sg13g2_decap_4
XFILLER_18_650 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1
+ VPWR VGND net2981 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2
+ net3104 i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2752 sg13g2_a221oi_1
XFILLER_33_686 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3060 net1336 net3066 net1322 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_mux2_1_A1
+ net1042 net568 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[380\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[380\]
+ net3126 i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2_sg13g2_a21o_1_X
+ net100 net3082 i_req_arb.data_i\[43\] i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y_sg13g2_inv_1_A
+ net94 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 VPWR VGND
+ sg13g2_inv_4
XFILLER_88_815 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2878
+ net2898 VPWR VGND sg13g2_nand2_1
XFILLER_29_904 VPWR VGND sg13g2_fill_2
XFILLER_101_168 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_A1
+ net1373 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net920 net2665 net2769 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1_Y
+ net2993 i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_nand2b_1_A_N_Y net3023 i_snitch.i_snitch_regfile.mem\[56\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_28_414 VPWR VGND sg13g2_fill_1
XFILLER_83_542 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3040
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_28_447 VPWR VGND sg13g2_fill_1
XFILLER_56_789 VPWR VGND sg13g2_fill_2
XFILLER_43_406 VPWR VGND sg13g2_fill_2
XFILLER_102_77 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_51_450 VPWR VGND sg13g2_fill_1
XFILLER_12_815 VPWR VGND sg13g2_fill_1
XFILLER_12_837 VPWR VGND sg13g2_fill_2
XFILLER_24_675 VPWR VGND sg13g2_decap_4
XFILLER_11_336 VPWR VGND sg13g2_decap_4
XFILLER_7_329 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[238\] clknet_leaf_88_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ net66 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2641 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_11_30 VPWR VGND sg13g2_fill_1
XFILLER_106_920 VPWR VGND sg13g2_decap_8
XFILLER_79_804 VPWR VGND sg13g2_fill_1
XFILLER_106_997 VPWR VGND sg13g2_decap_8
XFILLER_105_485 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2755 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_59_550 VPWR VGND sg13g2_decap_4
Xdata_pdata\[4\]_sg13g2_nor2_1_B net3161 data_pdata\[4\] data_pdata\[4\]_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_87_881 VPWR VGND sg13g2_decap_8
XFILLER_59_583 VPWR VGND sg13g2_decap_8
XFILLER_59_561 VPWR VGND sg13g2_fill_2
XFILLER_4_1004 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2650 VPWR VGND sg13g2_nand2_1
XFILLER_101_691 VPWR VGND sg13g2_decap_8
XFILLER_98_1011 VPWR VGND sg13g2_decap_8
XFILLER_74_520 VPWR VGND sg13g2_fill_1
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[0\]_sg13g2_dfrbpq_1_Q net3188 VGND VPWR net528 shift_reg_q\[0\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_27_491 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[453\]_sg13g2_nor3_1_A net1321 net2738 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_70_792 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net907 net2494 net1228 VPWR VGND sg13g2_a22oi_1
XFILLER_30_678 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net88 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
Xhold819 i_snitch.i_snitch_regfile.mem\[151\] VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold808 i_snitch.i_snitch_regfile.mem\[191\] VPWR VGND net840 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2860
+ net2657 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[76\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2354 net814 net2691 net2785 VPWR VGND sg13g2_a22oi_1
XFILLER_97_612 VPWR VGND sg13g2_fill_2
Xfanout3261 net3330 net3261 VPWR VGND sg13g2_buf_8
Xfanout3250 net3259 net3250 VPWR VGND sg13g2_buf_8
Xfanout3272 net3329 net3272 VPWR VGND sg13g2_buf_8
Xfanout3283 net3284 net3283 VPWR VGND sg13g2_buf_8
Xfanout2560 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y
+ net2560 VPWR VGND sg13g2_buf_8
Xfanout2571 net2575 net2571 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_69_358 VPWR VGND sg13g2_fill_2
Xi_snitch.gpr_waddr\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X net1389 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y i_snitch.gpr_waddr\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xfanout3294 net3300 net3294 VPWR VGND sg13g2_buf_8
Xfanout2582 net2583 net2582 VPWR VGND sg13g2_buf_1
XFILLER_97_689 VPWR VGND sg13g2_fill_1
XFILLER_96_155 VPWR VGND sg13g2_decap_4
Xfanout2593 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C_Y
+ net2593 VPWR VGND sg13g2_buf_8
XFILLER_65_542 VPWR VGND sg13g2_decap_8
XFILLER_38_756 VPWR VGND sg13g2_fill_1
XFILLER_65_575 VPWR VGND sg13g2_fill_1
XFILLER_65_564 VPWR VGND sg13g2_fill_2
XFILLER_93_895 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1_X
+ VPWR VGND sg13g2_and2_1
XFILLER_25_428 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[258\] clknet_leaf_109_clk sg13g2_dfrbpq_1
XFILLER_37_277 VPWR VGND sg13g2_fill_1
XFILLER_37_299 VPWR VGND sg13g2_fill_1
XFILLER_52_247 VPWR VGND sg13g2_decap_8
XFILLER_52_236 VPWR VGND sg13g2_decap_4
XFILLER_34_940 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_B
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ net2699 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.inst_addr_o\[22\] net2723 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ sg13g2_a21oi_1
Xtarget_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND target_sel_q_sg13g2_nand2b_1_A_N_Y sg13g2_nand2b_2
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y net2717
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2603 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_106_238 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[10\]_sg13g2_dfrbpq_1_Q net3239 VGND VPWR rsp_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[10\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2881
+ net2676 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2455
+ net2514 net2902 net2766 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2818 i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_103_956 VPWR VGND sg13g2_decap_8
XFILLER_102_477 VPWR VGND sg13g2_decap_4
XFILLER_88_689 VPWR VGND sg13g2_decap_4
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_69_870 VPWR VGND sg13g2_fill_1
XFILLER_29_745 VPWR VGND sg13g2_decap_8
XFILLER_84_884 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_decap_8
XFILLER_83_394 VPWR VGND sg13g2_decap_4
XFILLER_73_25 VPWR VGND sg13g2_fill_2
XFILLER_44_748 VPWR VGND sg13g2_decap_8
XFILLER_43_214 VPWR VGND sg13g2_decap_8
XFILLER_16_428 VPWR VGND sg13g2_fill_2
XFILLER_28_299 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2738
+ net2659 VPWR VGND sg13g2_nand2_1
XFILLER_24_450 VPWR VGND sg13g2_decap_4
XFILLER_25_973 VPWR VGND sg13g2_decap_4
XFILLER_40_910 VPWR VGND sg13g2_fill_2
XFILLER_106_1004 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[96\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[96\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2410 net872 net2904 net2869 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.inst_addr_o\[29\] net2524 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_12_678 VPWR VGND sg13g2_fill_1
XFILLER_7_137 VPWR VGND sg13g2_fill_1
XFILLER_7_115 VPWR VGND sg13g2_decap_4
XFILLER_11_188 VPWR VGND sg13g2_decap_4
Xi_snitch.consec_pc\[0\]_sg13g2_dfrbpq_1_Q net3260 VGND VPWR i_snitch.pc_d\[0\] i_snitch.consec_pc\[0\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_98_77 VPWR VGND sg13g2_decap_8
XFILLER_106_794 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_4_888 VPWR VGND sg13g2_fill_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_79_656 VPWR VGND sg13g2_decap_8
XFILLER_78_133 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[278\] clknet_leaf_65_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR net837 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_19_200 VPWR VGND sg13g2_fill_1
XFILLER_75_873 VPWR VGND sg13g2_fill_1
XFILLER_75_862 VPWR VGND sg13g2_fill_2
XFILLER_74_350 VPWR VGND sg13g2_fill_2
XFILLER_90_854 VPWR VGND sg13g2_decap_8
XFILLER_34_236 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2587 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[23\]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1 VGND VPWR i_snitch.inst_addr_o\[24\]
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[23\]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[23\]_sg13g2_mux2_1_A1_X sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[107\]
+ net2997 i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_43_770 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1_A2
+ VPWR VGND sg13g2_a21o_1
XFILLER_30_431 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[30\]_sg13g2_dfrbpq_1_Q net3244 VGND VPWR rsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[30\] clknet_leaf_39_clk sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net836 net715 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_30_497 VPWR VGND sg13g2_decap_4
Xhold627 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net659 sg13g2_dlygate4sd3_1
XFILLER_7_682 VPWR VGND sg13g2_fill_2
Xhold605 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\] VPWR
+ VGND net637 sg13g2_dlygate4sd3_1
Xhold616 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net648 sg13g2_dlygate4sd3_1
XFILLER_89_409 VPWR VGND sg13g2_fill_1
Xhold649 data_pdata\[7\] VPWR VGND net681 sg13g2_dlygate4sd3_1
Xhold638 i_snitch.i_snitch_regfile.mem\[283\] VPWR VGND net670 sg13g2_dlygate4sd3_1
XFILLER_98_976 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B VPWR
+ VGND sg13g2_and2_1
Xfanout3080 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1_X
+ net3080 VPWR VGND sg13g2_buf_8
Xfanout3091 net3093 net3091 VPWR VGND sg13g2_buf_8
XFILLER_97_464 VPWR VGND sg13g2_fill_2
XFILLER_85_615 VPWR VGND sg13g2_fill_1
Xhold1316 rsp_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1348
+ sg13g2_dlygate4sd3_1
Xi_snitch.sb_q\[14\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[14\] i_snitch.sb_q\[14\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
Xhold1305 i_snitch.i_snitch_regfile.mem\[357\] VPWR VGND net1337 sg13g2_dlygate4sd3_1
XFILLER_100_959 VPWR VGND sg13g2_decap_8
Xhold1349 rsp_data_q\[3\] VPWR VGND net1381 sg13g2_dlygate4sd3_1
XFILLER_66_840 VPWR VGND sg13g2_fill_2
Xdata_pdata\[12\]_sg13g2_nand2b_1_B data_pdata\[12\]_sg13g2_nand2b_1_B_Y data_pdata\[12\]
+ net3159 VPWR VGND sg13g2_nand2b_1
Xhold1338 i_snitch.i_snitch_regfile.mem\[133\] VPWR VGND net1370 sg13g2_dlygate4sd3_1
Xhold1327 i_snitch.i_snitch_regfile.mem\[259\] VPWR VGND net1359 sg13g2_dlygate4sd3_1
Xfanout2390 net2391 net2390 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[26\]_sg13g2_nand2_1_B i_snitch.pc_d\[26\]_sg13g2_nand2_1_B_Y i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[26\] VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2432 net2478 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_53_512 VPWR VGND sg13g2_fill_1
XFILLER_81_865 VPWR VGND sg13g2_decap_8
XFILLER_80_320 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ net2684 net2747 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_80_353 VPWR VGND sg13g2_fill_1
XFILLER_40_206 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[298\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ net2546 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ net2614 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[11\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net996 data_pdata\[11\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
XFILLER_1_825 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_89_965 VPWR VGND sg13g2_decap_8
XFILLER_102_252 VPWR VGND sg13g2_decap_8
XFILLER_76_604 VPWR VGND sg13g2_fill_1
XFILLER_0_379 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_1_1007 VPWR VGND sg13g2_decap_8
XFILLER_44_501 VPWR VGND sg13g2_fill_2
XFILLER_17_737 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2
+ net2633 VPWR i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y
+ VGND net2634 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2777 i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2906 net2430 i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q_D net2408
+ sg13g2_a221oi_1
XFILLER_71_375 VPWR VGND sg13g2_decap_8
XFILLER_44_589 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nor3_1_A net1288 net2782 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y
+ net2925 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ net3034 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A
+ VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
XFILLER_25_792 VPWR VGND sg13g2_fill_2
XFILLER_24_291 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C
+ net3141 VPWR VGND net3144 sg13g2_nand2b_2
XFILLER_12_475 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[117\] clknet_leaf_99_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[5\]
+ VGND net2293 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ VGND net2704 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xshift_reg_q\[16\]_sg13g2_dfrbpq_1_Q net3230 VGND VPWR net547 shift_reg_q\[16\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nor2b_1_B_N_Y
+ net3163 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[295\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_924 VPWR VGND sg13g2_decap_8
XFILLER_79_486 VPWR VGND sg13g2_fill_1
XFILLER_0_891 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2570 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ sg13g2_a21oi_1
XFILLER_75_692 VPWR VGND sg13g2_fill_2
XFILLER_63_843 VPWR VGND sg13g2_decap_8
XFILLER_22_206 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y
+ net2928 net51 net2848 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[64\]
+ i_snitch.i_snitch_regfile.mem\[96\] net3124 i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xdata_pdata\[31\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net859 data_pdata\[31\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2467 net2251 net2389 net1308 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VGND i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1 net3007 i_snitch.i_snitch_regfile.mem\[128\]
+ i_snitch.i_snitch_regfile.mem\[160\] i_snitch.i_snitch_regfile.mem\[192\] i_snitch.i_snitch_regfile.mem\[224\]
+ net2981 i_snitch.i_snitch_regfile.mem\[128\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_30_250 VPWR VGND sg13g2_fill_2
XFILLER_30_261 VPWR VGND sg13g2_fill_2
Xhold402 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\] VPWR
+ VGND net434 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[28\]_sg13g2_a22oi_1_A2_Y i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xhold435 i_snitch.i_snitch_regfile.mem\[377\] VPWR VGND net467 sg13g2_dlygate4sd3_1
Xhold413 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\] VPWR
+ VGND net445 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xhold424 i_snitch.i_snitch_regfile.mem\[306\] VPWR VGND net456 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[369\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2920
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y net2519 VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1
+ VGND i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xhold457 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net489 sg13g2_dlygate4sd3_1
Xhold468 cnt_q\[0\] VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold446 i_snitch.i_snitch_regfile.mem\[112\] VPWR VGND net478 sg13g2_dlygate4sd3_1
XFILLER_98_751 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y
+ net2539 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_nor2b_1
Xhold479 shift_reg_q\[23\] VPWR VGND net511 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_86_902 VPWR VGND sg13g2_decap_8
Xhold1102 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1134 sg13g2_dlygate4sd3_1
Xhold1124 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\] VPWR
+ VGND net1156 sg13g2_dlygate4sd3_1
Xhold1113 i_snitch.i_snitch_regfile.mem\[390\] VPWR VGND net1145 sg13g2_dlygate4sd3_1
XFILLER_100_756 VPWR VGND sg13g2_decap_8
XFILLER_86_979 VPWR VGND sg13g2_decap_8
Xhold1135 rsp_data_q\[24\] VPWR VGND net1167 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2379
+ sg13g2_o21ai_1
Xhold1146 i_snitch.i_snitch_regfile.mem\[178\] VPWR VGND net1178 sg13g2_dlygate4sd3_1
Xhold1157 i_snitch.i_snitch_regfile.mem\[501\] VPWR VGND net1189 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[137\] clknet_leaf_50_clk sg13g2_dfrbpq_1
Xhold1179 i_snitch.i_snitch_regfile.mem\[317\] VPWR VGND net1211 sg13g2_dlygate4sd3_1
XFILLER_26_501 VPWR VGND sg13g2_fill_1
Xhold1168 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\] VPWR
+ VGND net1200 sg13g2_dlygate4sd3_1
XFILLER_81_684 VPWR VGND sg13g2_decap_8
XFILLER_80_161 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_707 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ net2712 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_55_1020 VPWR VGND sg13g2_decap_8
XFILLER_6_928 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_nand2_1_B_Y
+ net3179 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\] VPWR
+ VGND sg13g2_nand2_1
Xshift_reg_q\[4\]_sg13g2_a22oi_1_A1 shift_reg_q\[4\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ net3057 net3047 net465 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[23\]_sg13g2_a21oi_1_A2 VGND VPWR net3160 data_pdata\[23\] data_pdata\[23\]_sg13g2_a21oi_1_A2_Y
+ net3152 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_nor3_1_A_Y net2454 net2765 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_dfrbpq_1_Q_D
+ net2909 sg13g2_a221oi_1
Xhold980 i_snitch.i_snitch_regfile.mem\[242\] VPWR VGND net1012 sg13g2_dlygate4sd3_1
Xhold991 i_snitch.i_snitch_regfile.mem\[243\] VPWR VGND net1023 sg13g2_dlygate4sd3_1
XFILLER_1_622 VPWR VGND sg13g2_decap_8
XFILLER_103_550 VPWR VGND sg13g2_fill_2
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_95_56 VPWR VGND sg13g2_decap_8
XFILLER_76_434 VPWR VGND sg13g2_decap_4
Xdata_pdata\[24\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2683 VPWR data_pdata\[24\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[24\]_sg13g2_nand2b_1_B_Y net3069 sg13g2_o21ai_1
XFILLER_0_176 VPWR VGND sg13g2_decap_8
XFILLER_1_699 VPWR VGND sg13g2_decap_8
XFILLER_92_927 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND net2706 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2546 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VGND net2585 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_85_990 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[433\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[433\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net792 net2663 net2864 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2958
+ i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2970
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_45_843 VPWR VGND sg13g2_fill_1
Xi_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.wake_up_q\[2\] clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_72_684 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_44_71 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_700 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2748 net2589 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2540 sg13g2_a21oi_1
XFILLER_5_32 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[157\] clknet_leaf_96_clk sg13g2_dfrbpq_1
XFILLER_95_710 VPWR VGND sg13g2_fill_2
XFILLER_86_209 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net960 net751 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_68_946 VPWR VGND sg13g2_fill_1
XFILLER_68_935 VPWR VGND sg13g2_decap_8
XFILLER_83_949 VPWR VGND sg13g2_decap_8
XFILLER_76_990 VPWR VGND sg13g2_decap_8
XFILLER_67_489 VPWR VGND sg13g2_decap_4
XFILLER_67_478 VPWR VGND sg13g2_fill_2
XFILLER_54_117 VPWR VGND sg13g2_fill_1
XFILLER_91_982 VPWR VGND sg13g2_decap_8
Xdata_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[6\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y
+ data_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y data_pdata\[30\]_sg13g2_a21oi_1_A2_Y
+ net3154 sg13g2_a21oi_2
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
XFILLER_50_345 VPWR VGND sg13g2_fill_1
XFILLER_50_334 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y
+ net2815 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_50_378 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_105_826 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_104_336 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2422 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_77_209 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_86_765 VPWR VGND sg13g2_fill_2
XFILLER_74_916 VPWR VGND sg13g2_fill_2
XFILLER_58_467 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2322
+ sg13g2_o21ai_1
XFILLER_105_77 VPWR VGND sg13g2_decap_8
XFILLER_100_575 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C_Y
+ VPWR VGND i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ sg13g2_nand3b_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_73_426 VPWR VGND sg13g2_fill_2
XFILLER_85_297 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B_sg13g2_o21ai_1_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B sg13g2_o21ai_1
XFILLER_54_651 VPWR VGND sg13g2_decap_4
XFILLER_26_364 VPWR VGND sg13g2_decap_8
XFILLER_82_993 VPWR VGND sg13g2_decap_8
XFILLER_81_470 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2757 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[177\] clknet_leaf_81_clk sg13g2_dfrbpq_1
XFILLER_10_732 VPWR VGND sg13g2_fill_2
XFILLER_6_725 VPWR VGND sg13g2_fill_2
XFILLER_5_213 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nor2b_1
XFILLER_6_758 VPWR VGND sg13g2_decap_8
XFILLER_100_0 VPWR VGND sg13g2_decap_8
Xfanout2912 data_pdata\[18\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2912 VPWR VGND
+ sg13g2_buf_8
Xfanout2901 net2902 net2901 VPWR VGND sg13g2_buf_8
Xfanout2923 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C
+ net2923 VPWR VGND sg13g2_buf_8
XFILLER_2_964 VPWR VGND sg13g2_decap_8
Xfanout2934 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2
+ net2934 VPWR VGND sg13g2_buf_8
Xfanout2945 net2946 net2945 VPWR VGND sg13g2_buf_8
Xfanout2967 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ net2967 VPWR VGND sg13g2_buf_8
XFILLER_49_401 VPWR VGND sg13g2_decap_8
Xfanout2978 net2979 net2978 VPWR VGND sg13g2_buf_8
Xfanout2989 net2995 net2989 VPWR VGND sg13g2_buf_8
Xfanout2956 net2960 net2956 VPWR VGND sg13g2_buf_8
XFILLER_65_916 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ VGND net2749 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
XFILLER_65_938 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_92_746 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_inv_1_Y
+ net2853 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2
+ VPWR VGND sg13g2_inv_4
XFILLER_64_459 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2417 sg13g2_a21oi_1
XFILLER_18_854 VPWR VGND sg13g2_fill_1
XFILLER_45_662 VPWR VGND sg13g2_fill_2
XFILLER_44_183 VPWR VGND sg13g2_fill_2
XFILLER_32_301 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[473\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[473\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net838 net2460 net2266 VPWR VGND sg13g2_a22oi_1
XFILLER_20_518 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0_X
+ net3096 net2931 i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q
+ net3188 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1
+ net90 VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y
+ VGND net2567 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2
+ sg13g2_o21ai_1
XFILLER_5_791 VPWR VGND sg13g2_fill_1
XFILLER_102_807 VPWR VGND sg13g2_decap_8
XFILLER_87_518 VPWR VGND sg13g2_fill_2
XFILLER_4_290 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2413
+ sg13g2_o21ai_1
XFILLER_95_551 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xor2_1
XFILLER_67_275 VPWR VGND sg13g2_fill_2
XFILLER_56_949 VPWR VGND sg13g2_decap_4
XFILLER_55_404 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2385
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2837 i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[364\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[364\] net2808 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[197\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[197\] clknet_leaf_118_clk sg13g2_dfrbpq_1
XFILLER_42_109 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[503\] clknet_leaf_67_clk sg13g2_dfrbpq_1
XFILLER_63_481 VPWR VGND sg13g2_fill_1
Xtarget_sel_q_sg13g2_nand2_1_B target_sel_q_sg13g2_nand2_1_B_Y net914 net1026 VPWR
+ VGND sg13g2_nand2_1
XFILLER_51_610 VPWR VGND sg13g2_fill_1
XFILLER_51_665 VPWR VGND sg13g2_decap_4
XFILLER_50_142 VPWR VGND sg13g2_fill_2
XFILLER_23_356 VPWR VGND sg13g2_decap_4
XFILLER_50_153 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[6\] net1133 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[331\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2399
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[45\] clknet_leaf_84_clk sg13g2_dfrbpq_1
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y net553
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C
+ i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2 VPWR VGND sg13g2_nor2_1
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_105_656 VPWR VGND sg13g2_decap_4
XFILLER_104_133 VPWR VGND sg13g2_decap_8
XFILLER_59_732 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2601 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_101_840 VPWR VGND sg13g2_decap_8
XFILLER_74_713 VPWR VGND sg13g2_decap_8
XFILLER_58_253 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[493\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2369 net1017 net2690 net2858 VPWR VGND sg13g2_a22oi_1
XFILLER_92_35 VPWR VGND sg13g2_decap_4
XFILLER_73_278 VPWR VGND sg13g2_fill_2
Xrebuffer91 net2608 net123 VPWR VGND sg13g2_buf_1
Xrebuffer80 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ net112 VPWR VGND sg13g2_buf_1
XFILLER_15_824 VPWR VGND sg13g2_decap_8
XFILLER_41_131 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q
+ net3191 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_10_540 VPWR VGND sg13g2_fill_1
XFILLER_6_533 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ net2575 VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1
+ VGND net2589 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_97_805 VPWR VGND sg13g2_decap_8
Xfanout2720 net2721 net2720 VPWR VGND sg13g2_buf_8
XFILLER_97_838 VPWR VGND sg13g2_decap_8
Xfanout2753 net2754 net2753 VPWR VGND sg13g2_buf_8
XFILLER_2_761 VPWR VGND sg13g2_decap_8
Xfanout2742 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2742 VPWR VGND sg13g2_buf_8
Xfanout2731 net2732 net2731 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D_sg13g2_or2_1_X
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y
+ net2566 sg13g2_or2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1
+ net2310 i_snitch.pc_d\[18\] i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
XFILLER_2_11 VPWR VGND sg13g2_decap_8
Xfanout2764 net2766 net2764 VPWR VGND sg13g2_buf_8
Xfanout2797 net2798 net2797 VPWR VGND sg13g2_buf_1
Xfanout2786 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X
+ net2786 VPWR VGND sg13g2_buf_8
Xfanout2775 net2776 net2775 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2666 net2780 net2318 net1246 VPWR VGND sg13g2_a22oi_1
XFILLER_2_88 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y
+ i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A VPWR
+ VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[65\] clknet_leaf_100_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2
+ net2305 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_B1
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2 VPWR
+ VGND i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_C1
+ net2761 net2965 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2852 sg13g2_a221oi_1
XFILLER_33_610 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y net556 VPWR i_snitch.sb_d\[12\] VGND net2293
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 net2515 VPWR VGND sg13g2_nand2_1
XFILLER_60_484 VPWR VGND sg13g2_fill_1
XFILLER_20_326 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[313\]
+ net3004 i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_a21oi_1_A1_Y net2977 sg13g2_a21oi_1
Xshift_reg_q\[21\]_sg13g2_nor2_1_A net483 net2728 shift_reg_q\[21\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_9_371 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_121_clk clknet_5_1__leaf_clk clknet_leaf_121_clk VPWR VGND sg13g2_buf_8
XFILLER_63_0 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y
+ net2561 net2601 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_0_709 VPWR VGND sg13g2_decap_8
XFILLER_102_648 VPWR VGND sg13g2_decap_8
XFILLER_101_147 VPWR VGND sg13g2_decap_8
Xcnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ net543 net500 VPWR VGND sg13g2_xnor2_1
XFILLER_68_562 VPWR VGND sg13g2_fill_2
XFILLER_56_702 VPWR VGND sg13g2_fill_2
XFILLER_83_532 VPWR VGND sg13g2_fill_2
XFILLER_83_565 VPWR VGND sg13g2_decap_8
XFILLER_83_587 VPWR VGND sg13g2_decap_8
XFILLER_71_749 VPWR VGND sg13g2_fill_2
XFILLER_102_56 VPWR VGND sg13g2_decap_8
XFILLER_62_27 VPWR VGND sg13g2_fill_2
Xdata_pdata\[6\]_sg13g2_dfrbpq_1_Q net3203 VGND VPWR net720 data_pdata\[6\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_24_687 VPWR VGND sg13g2_fill_1
XFILLER_11_315 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2889
+ net2693 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_112_clk clknet_5_16__leaf_clk clknet_leaf_112_clk VPWR VGND sg13g2_buf_8
XFILLER_20_871 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[100\]_sg13g2_nor3_1_A net1305 net2867 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2831 VPWR
+ i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a22oi_1_A1_Y sg13g2_o21ai_1
XFILLER_105_420 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2403 net949 net2691 net2796 VPWR VGND sg13g2_a22oi_1
Xcnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y net1 VPWR cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B1 sg13g2_o21ai_1
XFILLER_106_976 VPWR VGND sg13g2_decap_8
XFILLER_105_442 VPWR VGND sg13g2_fill_2
XFILLER_2_4 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[85\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_78_337 VPWR VGND sg13g2_decap_8
XFILLER_87_860 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]
+ net3176 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_2
XFILLER_19_404 VPWR VGND sg13g2_fill_1
XFILLER_100_191 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_440 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y
+ VGND sg13g2_inv_1
XFILLER_70_782 VPWR VGND sg13g2_fill_2
XFILLER_14_186 VPWR VGND sg13g2_fill_2
XFILLER_11_893 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2843
+ sg13g2_a221oi_1
Xclkbuf_leaf_103_clk clknet_5_19__leaf_clk clknet_leaf_103_clk VPWR VGND sg13g2_buf_8
Xhold809 i_snitch.i_snitch_regfile.mem\[41\] VPWR VGND net841 sg13g2_dlygate4sd3_1
Xdata_pdata\[1\]_sg13g2_mux2_1_A0 data_pdata\[1\] data_pdata\[9\] net3157 data_pdata\[1\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2597 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ net2587 sg13g2_a21oi_1
XFILLER_97_602 VPWR VGND sg13g2_fill_1
Xfanout3240 net3241 net3240 VPWR VGND sg13g2_buf_8
XFILLER_97_624 VPWR VGND sg13g2_decap_8
Xfanout3251 net3259 net3251 VPWR VGND sg13g2_buf_8
Xfanout3262 net3264 net3262 VPWR VGND sg13g2_buf_8
Xfanout3273 net3282 net3273 VPWR VGND sg13g2_buf_8
Xfanout2561 net2563 net2561 VPWR VGND sg13g2_buf_8
Xfanout2572 net2574 net2572 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ VGND net2749 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
Xfanout2550 net2553 net2550 VPWR VGND sg13g2_buf_8
XFILLER_85_808 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_Y
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y
+ sg13g2_nand4_1
Xfanout3284 net3287 net3284 VPWR VGND sg13g2_buf_8
Xfanout3295 net3300 net3295 VPWR VGND sg13g2_buf_8
Xfanout2594 net2595 net2594 VPWR VGND sg13g2_buf_8
Xfanout2583 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y
+ net2583 VPWR VGND sg13g2_buf_8
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
XFILLER_65_521 VPWR VGND sg13g2_decap_8
XFILLER_93_874 VPWR VGND sg13g2_decap_8
XFILLER_92_373 VPWR VGND sg13g2_fill_1
XFILLER_92_362 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2792
+ net2649 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
XFILLER_61_782 VPWR VGND sg13g2_fill_2
XFILLER_61_760 VPWR VGND sg13g2_decap_8
XFILLER_34_974 VPWR VGND sg13g2_fill_1
XFILLER_34_996 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2
+ net45 sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[352\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[352\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2398 net957 net2904 net2880 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2552 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2473 VPWR VGND sg13g2_nand2_1
XFILLER_106_217 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_103_935 VPWR VGND sg13g2_decap_8
XFILLER_88_624 VPWR VGND sg13g2_decap_4
XFILLER_87_101 VPWR VGND sg13g2_fill_1
XFILLER_0_539 VPWR VGND sg13g2_fill_2
XFILLER_87_178 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y
+ net2629 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_a22oi_1
XFILLER_68_370 VPWR VGND sg13g2_fill_1
XFILLER_84_863 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1167 net2497 net1374 VPWR VGND sg13g2_a22oi_1
XFILLER_56_576 VPWR VGND sg13g2_fill_1
XFILLER_25_930 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2562 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_24_484 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2478 net2460 i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2
+ VPWR VGND net2705 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1
+ net2547 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_3_300 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2581 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ net2577 sg13g2_a21oi_1
XFILLER_98_56 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q
+ net3230 VGND VPWR net636 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2876
+ net2653 VPWR VGND sg13g2_nand2_1
XFILLER_106_773 VPWR VGND sg13g2_decap_8
XFILLER_105_294 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_94_616 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1
+ net2722 i_snitch.inst_addr_o\[10\] i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
XFILLER_59_381 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B
+ net75 sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[372\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net985 net2672 net2882 VPWR VGND sg13g2_a22oi_1
XFILLER_75_885 VPWR VGND sg13g2_decap_8
XFILLER_74_373 VPWR VGND sg13g2_fill_2
XFILLER_47_587 VPWR VGND sg13g2_decap_4
XFILLER_47_93 VPWR VGND sg13g2_fill_1
XFILLER_35_716 VPWR VGND sg13g2_fill_1
XFILLER_50_708 VPWR VGND sg13g2_fill_1
XFILLER_72_1026 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2659 VPWR VGND sg13g2_nand2_1
XFILLER_31_933 VPWR VGND sg13g2_fill_2
XFILLER_31_955 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[373\]
+ net3119 i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_8_65 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2502 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2439 net2790 i_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[30\] net775 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xhold617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\] VPWR
+ VGND net649 sg13g2_dlygate4sd3_1
XFILLER_7_694 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[507\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2253 net2367 net1222 VPWR VGND sg13g2_a22oi_1
Xhold606 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net638 sg13g2_dlygate4sd3_1
Xhold639 i_snitch.i_snitch_regfile.mem\[286\] VPWR VGND net671 sg13g2_dlygate4sd3_1
Xhold628 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\] VPWR
+ VGND net660 sg13g2_dlygate4sd3_1
XFILLER_40_2 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VGND net2559 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_98_955 VPWR VGND sg13g2_decap_8
Xfanout3081 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1_X
+ net3081 VPWR VGND sg13g2_buf_8
Xfanout3070 i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_or2_1_A_X net3070 VPWR VGND
+ sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[402\] clknet_leaf_91_clk sg13g2_dfrbpq_1
Xfanout2380 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2380 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net1057 net2664 net2769 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1 VPWR VGND net3106 net2822
+ i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[61\]
+ i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1_Y net2827 sg13g2_a221oi_1
Xfanout3092 net3093 net3092 VPWR VGND sg13g2_buf_2
Xhold1306 i_snitch.i_snitch_regfile.mem\[228\] VPWR VGND net1338 sg13g2_dlygate4sd3_1
XFILLER_100_938 VPWR VGND sg13g2_decap_8
XFILLER_97_498 VPWR VGND sg13g2_fill_1
Xhold1317 rsp_data_q\[17\] VPWR VGND net1349 sg13g2_dlygate4sd3_1
Xhold1339 i_snitch.i_snitch_regfile.mem\[403\] VPWR VGND net1371 sg13g2_dlygate4sd3_1
Xhold1328 i_snitch.i_snitch_regfile.mem\[195\] VPWR VGND net1360 sg13g2_dlygate4sd3_1
Xfanout2391 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2391 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1
+ net806 net629 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_65_384 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VGND net2606 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_81_844 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_53_579 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2895
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_25_259 VPWR VGND sg13g2_fill_2
XFILLER_34_760 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ net69 VPWR VGND sg13g2_nand2_1
XFILLER_80_387 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2658 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\]_sg13g2_dfrbpq_1_Q
+ net3195 VGND VPWR net661 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
Xi_snitch.sb_q\[8\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.sb_d\[8\] i_snitch.sb_q\[8\]
+ clknet_leaf_106_clk sg13g2_dfrbpq_2
XFILLER_88_1022 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y net3116 sg13g2_o21ai_1
XFILLER_4_119 VPWR VGND sg13g2_decap_8
XFILLER_104_7 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[392\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net760 net2644 net3041 VPWR VGND sg13g2_a22oi_1
XFILLER_0_303 VPWR VGND sg13g2_fill_2
XFILLER_1_804 VPWR VGND sg13g2_decap_8
XFILLER_89_944 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A
+ net39 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor4_1
XFILLER_102_231 VPWR VGND sg13g2_decap_8
XFILLER_88_476 VPWR VGND sg13g2_fill_1
XFILLER_88_465 VPWR VGND sg13g2_decap_8
XFILLER_49_808 VPWR VGND sg13g2_decap_4
XFILLER_0_358 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2861
+ net2661 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2596 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_76_627 VPWR VGND sg13g2_decap_8
XFILLER_95_1015 VPWR VGND sg13g2_decap_8
XFILLER_57_896 VPWR VGND sg13g2_decap_4
XFILLER_57_885 VPWR VGND sg13g2_decap_8
XFILLER_16_215 VPWR VGND sg13g2_decap_8
XFILLER_17_716 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_fill_2
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_12_421 VPWR VGND sg13g2_fill_1
XFILLER_33_51 VPWR VGND sg13g2_fill_1
XFILLER_12_487 VPWR VGND sg13g2_decap_8
XFILLER_40_785 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y net2512
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2485 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2430 net657 i_snitch.i_snitch_regfile.mem\[290\]_sg13g2_dfrbpq_1_Q_D net2316
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[422\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_99_719 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[211\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net863 net2439 net2270 VPWR VGND sg13g2_a22oi_1
XFILLER_4_675 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2 net2831
+ VPWR i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_a21oi_1_A1_1_Y i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_4_697 VPWR VGND sg13g2_fill_1
XFILLER_95_903 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_and4_1_D
+ net3 net1122 net645 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C
+ VPWR VGND sg13g2_and4_1
XFILLER_0_870 VPWR VGND sg13g2_decap_8
XFILLER_94_468 VPWR VGND sg13g2_fill_1
XFILLER_94_457 VPWR VGND sg13g2_decap_8
XFILLER_75_682 VPWR VGND sg13g2_fill_2
Xstate_sg13g2_inv_1_A state_sg13g2_inv_1_A_Y state VPWR VGND sg13g2_inv_2
XFILLER_62_321 VPWR VGND sg13g2_decap_4
XFILLER_62_310 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_50_516 VPWR VGND sg13g2_fill_1
XFILLER_35_579 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_43_590 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[102\]
+ net2950 sg13g2_o21ai_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor3_2
Xhold403 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net435 sg13g2_dlygate4sd3_1
Xdata_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C i_snitch.i_snitch_lsu.metadata_q\[1\]
+ data_pdata\[20\]_sg13g2_mux2_1_A0_X data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y
+ VPWR VGND net3152 sg13g2_nand3b_1
Xhold436 shift_reg_q\[10\] VPWR VGND net468 sg13g2_dlygate4sd3_1
Xhold414 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold425 i_snitch.i_snitch_regfile.mem\[353\] VPWR VGND net457 sg13g2_dlygate4sd3_1
XFILLER_89_207 VPWR VGND sg13g2_decap_8
Xhold458 i_snitch.sb_q\[15\] VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold469 strb_reg_q\[0\] VPWR VGND net501 sg13g2_dlygate4sd3_1
Xhold447 shift_reg_q\[2\] VPWR VGND net479 sg13g2_dlygate4sd3_1
XFILLER_86_958 VPWR VGND sg13g2_decap_8
XFILLER_85_435 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2490 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X
+ sg13g2_o21ai_1
Xhold1114 i_snitch.i_snitch_regfile.mem\[434\] VPWR VGND net1146 sg13g2_dlygate4sd3_1
Xhold1103 i_snitch.i_snitch_regfile.mem\[166\] VPWR VGND net1135 sg13g2_dlygate4sd3_1
Xhold1125 rsp_data_q\[30\] VPWR VGND net1157 sg13g2_dlygate4sd3_1
Xhold1158 i_snitch.i_snitch_regfile.mem\[188\] VPWR VGND net1190 sg13g2_dlygate4sd3_1
Xhold1147 i_snitch.i_snitch_regfile.mem\[409\] VPWR VGND net1179 sg13g2_dlygate4sd3_1
Xhold1136 i_snitch.i_snitch_regfile.mem\[42\] VPWR VGND net1168 sg13g2_dlygate4sd3_1
XFILLER_39_863 VPWR VGND sg13g2_fill_1
XFILLER_94_980 VPWR VGND sg13g2_decap_8
Xhold1169 i_snitch.i_snitch_regfile.mem\[124\] VPWR VGND net1201 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_92_clk clknet_5_20__leaf_clk clknet_leaf_92_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2453 VPWR VGND sg13g2_nand2_1
XFILLER_38_384 VPWR VGND sg13g2_decap_4
XFILLER_38_395 VPWR VGND sg13g2_decap_8
XFILLER_53_365 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[442\] clknet_leaf_121_clk sg13g2_dfrbpq_1
XFILLER_26_579 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net962 net2451 net2267 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[231\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[231\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net1064 net2436 net2284 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2385
+ sg13g2_o21ai_1
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_22_785 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[196\]_sg13g2_nor3_1_A net1329 net2790 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[196\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_103_1019 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y
+ net2623 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[174\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1_sg13g2_inv_1_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1
+ i_snitch.sb_q\[12\] VGND sg13g2_inv_1
XFILLER_1_601 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C
+ VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B
+ sg13g2_nor4_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
Xhold970 i_snitch.i_snitch_regfile.mem\[173\] VPWR VGND net1002 sg13g2_dlygate4sd3_1
Xhold981 i_snitch.i_snitch_regfile.mem\[38\] VPWR VGND net1013 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B
+ net3035 net108 VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q
+ net3235 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
Xhold992 i_snitch.i_snitch_regfile.mem\[252\] VPWR VGND net1024 sg13g2_dlygate4sd3_1
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_1_678 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_95_35 VPWR VGND sg13g2_decap_8
XFILLER_92_906 VPWR VGND sg13g2_decap_8
XFILLER_76_446 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2728 shift_reg_q\[13\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[9\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[9\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_91_427 VPWR VGND sg13g2_decap_8
XFILLER_63_107 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ VGND net2600 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_57_693 VPWR VGND sg13g2_fill_1
XFILLER_29_384 VPWR VGND sg13g2_decap_8
XFILLER_29_395 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_83_clk clknet_5_23__leaf_clk clknet_leaf_83_clk VPWR VGND sg13g2_buf_8
XFILLER_71_151 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[23\]_sg13g2_dfrbpq_1_Q net3237 VGND VPWR rsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[23\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_44_94 VPWR VGND sg13g2_decap_4
XFILLER_44_83 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_734 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ sg13g2_nand2b_2
XFILLER_5_11 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_5_984 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[410\]
+ i_snitch.i_snitch_regfile.mem\[442\] i_snitch.i_snitch_regfile.mem\[474\] i_snitch.i_snitch_regfile.mem\[506\]
+ net3099 i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_99_538 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C
+ VGND net2541 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_95_700 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[462\] clknet_leaf_82_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_A1
+ net1197 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[251\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net782 net2436 net2252 VPWR VGND sg13g2_a22oi_1
XFILLER_83_928 VPWR VGND sg13g2_decap_8
Xuo_out_sg13g2_buf_1_X req_data_valid net17 VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_74_clk clknet_5_25__leaf_clk clknet_leaf_74_clk VPWR VGND sg13g2_buf_8
XFILLER_91_961 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_36_888 VPWR VGND sg13g2_fill_2
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
XFILLER_90_482 VPWR VGND sg13g2_decap_8
XFILLER_51_825 VPWR VGND sg13g2_fill_2
XFILLER_93_0 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B_sg13g2_a221oi_1_C1
+ VPWR VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2421 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[458\]_sg13g2_o21ai_1_A1 net2962 VPWR i_snitch.i_snitch_regfile.mem\[458\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[458\] i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[480\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y net2957
+ i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2969
+ i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2627 net2853 net3084
+ VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q
+ net3188 VGND VPWR net602 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_105_805 VPWR VGND sg13g2_decap_8
XFILLER_85_1025 VPWR VGND sg13g2_decap_4
XFILLER_104_315 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_fill_2
XFILLER_98_593 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2322
+ sg13g2_o21ai_1
XFILLER_105_56 VPWR VGND sg13g2_decap_8
XFILLER_86_777 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B_Y VPWR
+ VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ sg13g2_nand3b_1
XFILLER_73_449 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_65_clk clknet_5_25__leaf_clk clknet_leaf_65_clk VPWR VGND sg13g2_buf_8
XFILLER_26_310 VPWR VGND sg13g2_fill_1
XFILLER_82_972 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_decap_4
XFILLER_27_866 VPWR VGND sg13g2_fill_1
XFILLER_27_888 VPWR VGND sg13g2_fill_1
XFILLER_92_1018 VPWR VGND sg13g2_decap_8
XFILLER_81_493 VPWR VGND sg13g2_decap_4
XFILLER_26_376 VPWR VGND sg13g2_decap_4
XFILLER_42_847 VPWR VGND sg13g2_fill_1
XFILLER_41_379 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0 net3123 i_snitch.i_snitch_regfile.mem\[136\]
+ i_snitch.i_snitch_regfile.mem\[168\] i_snitch.i_snitch_regfile.mem\[200\] i_snitch.i_snitch_regfile.mem\[232\]
+ net3113 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_10_766 VPWR VGND sg13g2_decap_4
XFILLER_5_203 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[482\] clknet_leaf_109_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D_sg13g2_nor2_1_Y
+ net3085 net3083 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_nor2_1
Xdata_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[0\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y
+ data_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y data_pdata\[24\]_sg13g2_a21oi_1_A2_Y
+ net3152 sg13g2_a21oi_2
Xdata_pdata\[25\]_sg13g2_nand2b_1_B data_pdata\[25\]_sg13g2_nand2b_1_B_Y data_pdata\[25\]
+ VPWR VGND net3155 sg13g2_nand2b_2
Xi_snitch.i_snitch_regfile.mem\[271\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2326 net1030 net2677 net2894 VPWR VGND sg13g2_a22oi_1
XFILLER_5_258 VPWR VGND sg13g2_fill_2
XFILLER_30_52 VPWR VGND sg13g2_fill_2
XFILLER_2_943 VPWR VGND sg13g2_decap_8
Xfanout2902 data_pdata\[25\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2902 VPWR
+ VGND sg13g2_buf_8
XFILLER_96_519 VPWR VGND sg13g2_decap_4
Xfanout2924 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2
+ net2924 VPWR VGND sg13g2_buf_8
Xfanout2913 net2914 net2913 VPWR VGND sg13g2_buf_8
Xfanout2946 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net2946 VPWR VGND sg13g2_buf_8
Xfanout2935 net2939 net2935 VPWR VGND sg13g2_buf_8
XFILLER_104_893 VPWR VGND sg13g2_decap_8
Xfanout2957 net2960 net2957 VPWR VGND sg13g2_buf_2
Xfanout2968 net2969 net2968 VPWR VGND sg13g2_buf_8
XFILLER_7_1025 VPWR VGND sg13g2_decap_4
Xfanout2979 net2996 net2979 VPWR VGND sg13g2_buf_8
XFILLER_103_392 VPWR VGND sg13g2_decap_8
XFILLER_77_744 VPWR VGND sg13g2_fill_2
XFILLER_76_221 VPWR VGND sg13g2_fill_1
XFILLER_49_435 VPWR VGND sg13g2_fill_2
XFILLER_91_202 VPWR VGND sg13g2_fill_2
XFILLER_49_468 VPWR VGND sg13g2_decap_8
XFILLER_36_107 VPWR VGND sg13g2_fill_2
XFILLER_92_769 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_56_clk clknet_5_31__leaf_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2861 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2
+ net2505 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_72_471 VPWR VGND sg13g2_decap_4
XFILLER_60_600 VPWR VGND sg13g2_fill_2
Xdata_pdata\[24\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net928 data_pdata\[24\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_2
XFILLER_60_633 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[406\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2391 net1100 net2652 net3042 VPWR VGND sg13g2_a22oi_1
XFILLER_32_324 VPWR VGND sg13g2_fill_1
XFILLER_60_688 VPWR VGND sg13g2_decap_8
XFILLER_32_379 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[301\] clknet_leaf_85_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B
+ net3016 net2997 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y
+ net1332 i_req_arb.gen_arbiter.req_d\[1\] i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2818 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_99_379 VPWR VGND sg13g2_decap_8
XFILLER_45_1020 VPWR VGND sg13g2_decap_8
XFILLER_101_329 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[75\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[75\]
+ i_snitch.i_snitch_regfile.mem\[107\] net3136 i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2840
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[1\] net954 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2 i_snitch.pc_d\[12\]_sg13g2_mux2_1_A1_A0
+ VPWR VGND sg13g2_and2_1
XFILLER_67_254 VPWR VGND sg13g2_fill_1
XFILLER_95_596 VPWR VGND sg13g2_fill_2
XFILLER_83_758 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2363
+ sg13g2_o21ai_1
XFILLER_49_991 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2_sg13g2_nand3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2535 i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_A i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2
+ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_47_clk clknet_5_13__leaf_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
XFILLER_23_302 VPWR VGND sg13g2_decap_4
XFILLER_24_825 VPWR VGND sg13g2_decap_4
XFILLER_35_173 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2696 net2541 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[308\] net3020 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_nand3_1
Xdata_pdata\[16\]_sg13g2_a21oi_1_A2 VGND VPWR net3159 data_pdata\[16\] data_pdata\[16\]_sg13g2_a21oi_1_A2_Y
+ net3152 sg13g2_a21oi_1
XFILLER_3_707 VPWR VGND sg13g2_decap_8
XFILLER_105_635 VPWR VGND sg13g2_fill_1
XFILLER_104_112 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y_sg13g2_nand3_1_A
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_C
+ VPWR VGND sg13g2_nand3_1
XFILLER_78_519 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[292\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[292\]
+ net3007 i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_a21oi_1_A1_Y net2980 sg13g2_a21oi_1
XFILLER_104_189 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[2\]_sg13g2_nor2_1_A net479 net2731 shift_reg_q\[2\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[120\]
+ net2952 i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_59_744 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[426\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2465 net2283 net2381 net1185 VPWR VGND sg13g2_a22oi_1
XFILLER_47_917 VPWR VGND sg13g2_fill_2
XFILLER_101_896 VPWR VGND sg13g2_decap_8
XFILLER_100_373 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_38_clk clknet_5_10__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_92_14 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[321\] clknet_leaf_76_clk sg13g2_dfrbpq_1
Xrebuffer70 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C
+ net102 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y VPWR
+ VGND sg13g2_nand2_2
Xrebuffer81 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ net113 VPWR VGND sg13g2_buf_1
XFILLER_15_814 VPWR VGND sg13g2_fill_2
XFILLER_26_151 VPWR VGND sg13g2_fill_1
XFILLER_27_696 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2570 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xrebuffer92 net3128 net124 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2411 net911 net2688 net2870 VPWR VGND sg13g2_a22oi_1
XFILLER_30_806 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ net2853 VPWR VGND sg13g2_nand2_1
XFILLER_10_574 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B_sg13g2_nor2_1_Y
+ i_snitch.inst_addr_o\[12\] net2527 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2424 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[161\]_sg13g2_nand2_1_A_1 i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_nand2_1_A_1_Y
+ i_snitch.i_snitch_regfile.mem\[161\] net2826 VPWR VGND sg13g2_nand2_1
XFILLER_97_817 VPWR VGND sg13g2_decap_8
Xfanout2710 net2711 net2710 VPWR VGND sg13g2_buf_1
Xfanout2721 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X
+ net2721 VPWR VGND sg13g2_buf_8
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1
+ net540 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
XFILLER_2_740 VPWR VGND sg13g2_decap_8
Xfanout2754 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y
+ net2754 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2321
+ sg13g2_o21ai_1
Xfanout2743 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ net2743 VPWR VGND sg13g2_buf_8
XFILLER_1_261 VPWR VGND sg13g2_fill_2
Xfanout2732 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y net2732
+ VPWR VGND sg13g2_buf_8
Xfanout2765 net2766 net2765 VPWR VGND sg13g2_buf_1
Xfanout2776 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1_X
+ net2776 VPWR VGND sg13g2_buf_8
Xfanout2787 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X
+ net2787 VPWR VGND sg13g2_buf_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
Xfanout2798 net2799 net2798 VPWR VGND sg13g2_buf_8
XFILLER_37_416 VPWR VGND sg13g2_fill_1
XFILLER_37_438 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C
+ net2548 VGND sg13g2_inv_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y net2717
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_29_clk clknet_5_8__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_64_246 VPWR VGND sg13g2_fill_1
XFILLER_52_408 VPWR VGND sg13g2_decap_8
XFILLER_46_972 VPWR VGND sg13g2_fill_2
XFILLER_46_961 VPWR VGND sg13g2_fill_2
XFILLER_92_599 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ VPWR VGND sg13g2_and2_1
XFILLER_75_1013 VPWR VGND sg13g2_decap_8
XFILLER_61_942 VPWR VGND sg13g2_decap_8
XFILLER_45_493 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]
+ net3179 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B_sg13g2_and3_1_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B
+ net3033 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ VPWR VGND sg13g2_and3_2
Xheichips25_snitch_wrapper_30 VPWR VGND uio_oe[2] sg13g2_tiehi
XFILLER_33_677 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2684 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_891 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ net1236 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
XFILLER_102_627 VPWR VGND sg13g2_fill_2
XFILLER_102_616 VPWR VGND sg13g2_fill_2
XFILLER_82_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q net3264 VGND VPWR i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[341\] clknet_leaf_113_clk sg13g2_dfrbpq_1
XFILLER_101_126 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_96_894 VPWR VGND sg13g2_decap_8
XFILLER_68_585 VPWR VGND sg13g2_fill_1
XFILLER_56_747 VPWR VGND sg13g2_decap_8
XFILLER_55_213 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[447\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[447\]
+ net3009 i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_a21oi_1_A1_Y net2983 sg13g2_a21oi_1
XFILLER_102_35 VPWR VGND sg13g2_decap_8
XFILLER_71_739 VPWR VGND sg13g2_decap_4
XFILLER_52_942 VPWR VGND sg13g2_decap_8
XFILLER_24_644 VPWR VGND sg13g2_decap_4
XFILLER_36_482 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2341
+ sg13g2_o21ai_1
XFILLER_12_839 VPWR VGND sg13g2_fill_1
XFILLER_23_176 VPWR VGND sg13g2_decap_4
XFILLER_7_309 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2640 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_11_21 VPWR VGND sg13g2_decap_8
XFILLER_106_955 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2706 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_93_319 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nand2b_1
Xdata_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A
+ VPWR data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y
+ data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VGND
+ sg13g2_inv_1
XFILLER_100_170 VPWR VGND sg13g2_decap_8
XFILLER_86_360 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_19_416 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B
+ net2499 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_961 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VGND net2588 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_74_588 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y net3163
+ net2487 i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 VPWR VGND
+ sg13g2_nor2_1
XFILLER_27_460 VPWR VGND sg13g2_fill_1
XFILLER_28_972 VPWR VGND sg13g2_fill_1
XFILLER_61_249 VPWR VGND sg13g2_decap_4
XFILLER_55_791 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[466\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net1123 net2461 net2273 VPWR VGND sg13g2_a22oi_1
XFILLER_42_452 VPWR VGND sg13g2_fill_2
XFILLER_11_850 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2605 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[361\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_10_371 VPWR VGND sg13g2_fill_2
XFILLER_10_360 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2463 net2860 i_snitch.i_snitch_regfile.mem\[419\]_sg13g2_dfrbpq_1_Q_D net2909
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ net2577 VPWR VGND sg13g2_a22oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D_sg13g2_or2_1_X
+ VGND VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ net3141 sg13g2_or2_1
Xdata_pdata\[1\]_sg13g2_mux2_1_A1 rsp_data_q\[1\] net734 net3048 data_pdata\[1\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xshift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ VPWR shift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 VGND net3172 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net853 net2651 net2888 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xfanout3230 net3232 net3230 VPWR VGND sg13g2_buf_8
Xfanout3241 net3249 net3241 VPWR VGND sg13g2_buf_8
XFILLER_69_316 VPWR VGND sg13g2_decap_4
Xfanout3252 net3253 net3252 VPWR VGND sg13g2_buf_8
Xfanout3263 net3264 net3263 VPWR VGND sg13g2_buf_8
Xfanout3274 net3282 net3274 VPWR VGND sg13g2_buf_8
Xfanout2562 net88 net2562 VPWR VGND sg13g2_buf_1
Xfanout2540 net2541 net2540 VPWR VGND sg13g2_buf_8
Xfanout2551 net2552 net2551 VPWR VGND sg13g2_buf_8
Xfanout3285 net3287 net3285 VPWR VGND sg13g2_buf_8
Xfanout3296 net3300 net3296 VPWR VGND sg13g2_buf_8
Xfanout2595 net2598 net2595 VPWR VGND sg13g2_buf_1
Xfanout2584 net2585 net2584 VPWR VGND sg13g2_buf_8
Xfanout2573 net2574 net2573 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1
+ net2722 i_snitch.inst_addr_o\[24\] i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_93_853 VPWR VGND sg13g2_decap_8
XFILLER_92_352 VPWR VGND sg13g2_fill_2
XFILLER_92_341 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[357\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[357\] net2801 sg13g2_o21ai_1
XFILLER_37_235 VPWR VGND sg13g2_decap_8
XFILLER_25_408 VPWR VGND sg13g2_fill_1
XFILLER_25_419 VPWR VGND sg13g2_decap_8
XFILLER_80_558 VPWR VGND sg13g2_fill_1
XFILLER_33_441 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.inst_addr_o\[21\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[21\]
+ i_snitch.inst_addr_o\[21\] clknet_leaf_58_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q net3280 VGND VPWR i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[38\] clknet_leaf_76_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xclkbuf_leaf_9_clk clknet_5_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_103_914 VPWR VGND sg13g2_decap_8
XFILLER_88_603 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_88_658 VPWR VGND sg13g2_decap_8
Xdata_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2 data_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ net3070 net2714 data_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 net2517 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ net2758 VPWR VGND sg13g2_a22oi_1
XFILLER_69_894 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[486\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2369 net878 net2900 net2858 VPWR VGND sg13g2_a22oi_1
XFILLER_84_842 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2934 i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_246 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ net85 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[381\] clknet_leaf_95_clk sg13g2_dfrbpq_1
XFILLER_71_569 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q
+ net3228 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_12_603 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[170\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[170\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2282 net2344 net1192
+ VPWR VGND sg13g2_a22oi_1
XFILLER_40_912 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y VGND
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ sg13g2_a21oi_1
XFILLER_40_945 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[487\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[487\]
+ net3117 i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_a21oi_1_A1_Y net2940 sg13g2_a21oi_1
XFILLER_7_128 VPWR VGND sg13g2_decap_8
XFILLER_11_157 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ net2578 VPWR VGND sg13g2_a22oi_1
XFILLER_98_35 VPWR VGND sg13g2_decap_8
XFILLER_106_752 VPWR VGND sg13g2_decap_8
XFILLER_106_741 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_mux2_1_X
+ net47 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net2709 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_4_846 VPWR VGND sg13g2_decap_8
XFILLER_79_625 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[377\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[377\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[377\] net2800 sg13g2_o21ai_1
XFILLER_105_273 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_2
XFILLER_79_669 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[305\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2663 net2781 net2319 net1266 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2704 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_75_864 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[58\] clknet_leaf_113_clk sg13g2_dfrbpq_1
XFILLER_19_235 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X
+ net2486 i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q_D i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[200\] clknet_leaf_73_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[478\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B i_snitch.consec_pc\[0\] i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_90_889 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_15_430 VPWR VGND sg13g2_fill_1
XFILLER_16_964 VPWR VGND sg13g2_decap_8
XFILLER_97_7 VPWR VGND sg13g2_decap_8
XFILLER_15_485 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_A1
+ net2303 i_snitch.pc_d\[29\] i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_nor3_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A_C
+ VPWR VGND sg13g2_nor3_1
XFILLER_7_640 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold607 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\] VPWR
+ VGND net639 sg13g2_dlygate4sd3_1
Xhold618 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net650 sg13g2_dlygate4sd3_1
XFILLER_7_684 VPWR VGND sg13g2_fill_1
XFILLER_7_673 VPWR VGND sg13g2_fill_2
Xhold629 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[42\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net661 sg13g2_dlygate4sd3_1
XFILLER_98_934 VPWR VGND sg13g2_decap_8
XFILLER_97_433 VPWR VGND sg13g2_fill_1
Xfanout3060 net3061 net3060 VPWR VGND sg13g2_buf_8
Xfanout3082 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1_X
+ net3082 VPWR VGND sg13g2_buf_8
Xfanout3071 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ net3071 VPWR VGND sg13g2_buf_8
XFILLER_100_917 VPWR VGND sg13g2_decap_8
XFILLER_97_466 VPWR VGND sg13g2_fill_1
Xfanout3093 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_X
+ net3093 VPWR VGND sg13g2_buf_8
Xfanout2370 net2371 net2370 VPWR VGND sg13g2_buf_8
Xhold1307 i_snitch.i_snitch_regfile.mem\[418\] VPWR VGND net1339 sg13g2_dlygate4sd3_1
Xdata_pdata\[1\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B net3149 data_pdata\[1\]_sg13g2_mux2_1_A0_X
+ data_pdata\[1\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
XFILLER_78_680 VPWR VGND sg13g2_decap_4
Xhold1318 rsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1350
+ sg13g2_dlygate4sd3_1
Xhold1329 i_req_arb.data_i\[41\] VPWR VGND net1361 sg13g2_dlygate4sd3_1
Xfanout2392 net2393 net2392 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[190\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y net2244 net2344 net1244
+ VPWR VGND sg13g2_a22oi_1
Xfanout2381 net2383 net2381 VPWR VGND sg13g2_buf_8
XFILLER_19_0 VPWR VGND sg13g2_fill_2
XFILLER_92_160 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_nor2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A VPWR VGND sg13g2_nor2_2
XFILLER_66_886 VPWR VGND sg13g2_decap_4
XFILLER_38_566 VPWR VGND sg13g2_fill_2
XFILLER_53_547 VPWR VGND sg13g2_fill_1
XFILLER_19_780 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1365 net2491 net1258 VPWR VGND sg13g2_a22oi_1
XFILLER_21_400 VPWR VGND sg13g2_fill_1
XFILLER_22_945 VPWR VGND sg13g2_decap_8
XFILLER_21_444 VPWR VGND sg13g2_fill_2
XFILLER_88_1001 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2638 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[155\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_A1 net2524 VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1
+ net2590 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_nor2_1_B
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_89_923 VPWR VGND sg13g2_decap_8
XFILLER_88_400 VPWR VGND sg13g2_decap_8
Xdata_pdata\[8\]_sg13g2_mux2_1_A1 rsp_data_q\[8\] net1147 net3051 data_pdata\[8\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[78\] clknet_leaf_83_clk sg13g2_dfrbpq_1
XFILLER_102_210 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[220\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net3162 net2486 i_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_103_788 VPWR VGND sg13g2_decap_8
XFILLER_102_287 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1_Y
+ VGND net2709 i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_84_683 VPWR VGND sg13g2_decap_8
XFILLER_84_661 VPWR VGND sg13g2_fill_2
XFILLER_44_503 VPWR VGND sg13g2_fill_1
XFILLER_17_739 VPWR VGND sg13g2_fill_1
XFILLER_44_569 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[167\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2771
+ net2897 VPWR VGND sg13g2_nand2_1
XFILLER_13_967 VPWR VGND sg13g2_decap_8
XFILLER_8_426 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2789
+ net2655 VPWR VGND sg13g2_nand2_1
XFILLER_8_448 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_Y
+ net2490 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2b_1
XFILLER_4_654 VPWR VGND sg13g2_decap_8
XFILLER_106_593 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_39_308 VPWR VGND sg13g2_decap_4
XFILLER_95_959 VPWR VGND sg13g2_decap_8
XFILLER_94_403 VPWR VGND sg13g2_fill_2
XFILLER_66_116 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ net2696 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y net2718
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_63_834 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y
+ net67 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nor2_1
XFILLER_90_686 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net781 net2472 net2267 VPWR VGND sg13g2_a22oi_1
XFILLER_16_772 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[98\] clknet_leaf_108_clk sg13g2_dfrbpq_1
XFILLER_30_252 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A_Y net2843 i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q net3289 VGND VPWR i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[240\] clknet_leaf_89_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B
+ net2958 i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xhold404 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\] VPWR
+ VGND net436 sg13g2_dlygate4sd3_1
Xhold426 i_snitch.i_snitch_regfile.mem\[65\] VPWR VGND net458 sg13g2_dlygate4sd3_1
Xhold415 i_snitch.i_snitch_regfile.mem\[481\] VPWR VGND net447 sg13g2_dlygate4sd3_1
Xhold459 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1 VPWR VGND net491 sg13g2_dlygate4sd3_1
Xhold437 shift_reg_q\[10\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net469 sg13g2_dlygate4sd3_1
Xhold448 shift_reg_q\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net480 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2440 VPWR VGND sg13g2_nand2_1
XFILLER_97_263 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[4\]_sg13g2_dfrbpq_1_Q net3241 VGND VPWR rsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[4\] clknet_leaf_38_clk sg13g2_dfrbpq_2
XFILLER_86_937 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y
+ i_snitch.inst_addr_o\[30\] i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1 VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2735 shift_reg_q\[24\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[20\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[20\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold1115 data_pdata\[8\] VPWR VGND net1147 sg13g2_dlygate4sd3_1
Xhold1104 i_snitch.i_snitch_regfile.mem\[506\] VPWR VGND net1136 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ net3098 i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ net2918 sg13g2_a221oi_1
XFILLER_100_747 VPWR VGND sg13g2_decap_4
Xhold1126 rsp_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1158
+ sg13g2_dlygate4sd3_1
Xhold1137 rsp_data_q\[22\] VPWR VGND net1169 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2872
+ net2657 VPWR VGND sg13g2_nand2_1
Xhold1148 i_snitch.i_snitch_regfile.mem\[125\] VPWR VGND net1180 sg13g2_dlygate4sd3_1
XFILLER_39_831 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A
+ VGND net2541 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xhold1159 i_snitch.i_snitch_regfile.mem\[376\] VPWR VGND net1191 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ VPWR i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y
+ VGND net2959 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2
+ sg13g2_o21ai_1
XFILLER_26_536 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[344\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2379
+ sg13g2_o21ai_1
XFILLER_41_528 VPWR VGND sg13g2_decap_4
XFILLER_80_196 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\] net616 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q VPWR VGND
+ sg13g2_nand2_1
XFILLER_70_39 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X
+ net2810 net2818 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y
+ VPWR VGND sg13g2_nor4_1
XFILLER_10_948 VPWR VGND sg13g2_fill_2
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1_sg13g2_nand2_1_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR net575 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ net64 net2519 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1 VPWR VGND sg13g2_nand3_1
XFILLER_89_742 VPWR VGND sg13g2_fill_1
Xhold971 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] VPWR
+ VGND net1003 sg13g2_dlygate4sd3_1
Xhold960 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net992 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nand4_1_A i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_Y i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y
+ i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_C VPWR VGND i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A_Y
+ sg13g2_nand4_1
XFILLER_0_112 VPWR VGND sg13g2_decap_8
Xhold982 i_snitch.i_snitch_regfile.mem\[365\] VPWR VGND net1014 sg13g2_dlygate4sd3_1
XFILLER_103_530 VPWR VGND sg13g2_decap_8
XFILLER_95_14 VPWR VGND sg13g2_decap_8
Xhold993 i_snitch.i_snitch_regfile.mem\[491\] VPWR VGND net1025 sg13g2_dlygate4sd3_1
XFILLER_1_657 VPWR VGND sg13g2_decap_8
XFILLER_76_425 VPWR VGND sg13g2_fill_2
XFILLER_76_414 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net1014 net2689 net2881 VPWR VGND sg13g2_a22oi_1
XFILLER_91_417 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2695 net2599 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q net3250 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\] clknet_leaf_19_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2638 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q net3220 VGND VPWR i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[260\] clknet_leaf_107_clk sg13g2_dfrbpq_1
XFILLER_72_653 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ net3034 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y
+ VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
XFILLER_72_686 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_32_528 VPWR VGND sg13g2_fill_1
XFILLER_9_702 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 net2833
+ VPWR i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2817 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[366\]
+ net3130 i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_a21oi_1_A1_Y net2943 sg13g2_a21oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y
+ net2567 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_60_50 VPWR VGND sg13g2_decap_4
XFILLER_9_779 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[371\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2660 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2662 VPWR VGND sg13g2_nand2_1
XFILLER_99_528 VPWR VGND sg13g2_decap_4
XFILLER_5_963 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0_X
+ net2938 net2931 i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_95_745 VPWR VGND sg13g2_decap_8
XFILLER_83_907 VPWR VGND sg13g2_decap_8
XFILLER_48_661 VPWR VGND sg13g2_fill_2
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_94_299 VPWR VGND sg13g2_fill_1
XFILLER_91_940 VPWR VGND sg13g2_decap_8
XFILLER_78_1022 VPWR VGND sg13g2_decap_8
XFILLER_36_823 VPWR VGND sg13g2_fill_1
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_62_174 VPWR VGND sg13g2_decap_4
XFILLER_50_303 VPWR VGND sg13g2_decap_4
XFILLER_16_580 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR net437 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_86_0 VPWR VGND sg13g2_decap_8
XFILLER_31_561 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1157 net2495 net1181 VPWR VGND sg13g2_a22oi_1
XFILLER_85_1004 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ VGND VPWR net2848 sg13g2_nor4_2
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D
+ VGND net2610 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q net3315 VGND VPWR i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[280\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_98_561 VPWR VGND sg13g2_fill_2
XFILLER_86_734 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
XFILLER_105_35 VPWR VGND sg13g2_decap_8
XFILLER_86_767 VPWR VGND sg13g2_fill_1
XFILLER_86_745 VPWR VGND sg13g2_decap_4
XFILLER_74_918 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_85_288 VPWR VGND sg13g2_fill_2
XFILLER_73_428 VPWR VGND sg13g2_fill_1
XFILLER_82_951 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
XFILLER_81_461 VPWR VGND sg13g2_decap_8
XFILLER_26_399 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[276\]_sg13g2_o21ai_1_A1 net2937 VPWR i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[276\] net2814 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[415\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_10_734 VPWR VGND sg13g2_fill_1
XFILLER_6_727 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[204\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[204\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net926 net2692 net2791 VPWR VGND sg13g2_a22oi_1
XFILLER_6_749 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net458 net2353 VPWR VGND sg13g2_nand2_1
Xfanout2903 data_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2903 VPWR
+ VGND sg13g2_buf_8
XFILLER_2_922 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2415 sg13g2_a21oi_1
Xhold790 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\] VPWR
+ VGND net822 sg13g2_dlygate4sd3_1
Xfanout2925 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ net2925 VPWR VGND sg13g2_buf_8
Xfanout2914 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y net2914 VPWR
+ VGND sg13g2_buf_8
Xfanout2936 net2938 net2936 VPWR VGND sg13g2_buf_8
XFILLER_104_872 VPWR VGND sg13g2_decap_8
XFILLER_89_572 VPWR VGND sg13g2_decap_8
Xfanout2969 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2969 VPWR VGND sg13g2_buf_8
XFILLER_7_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_999 VPWR VGND sg13g2_decap_8
Xfanout2958 net2960 net2958 VPWR VGND sg13g2_buf_8
Xfanout2947 net2949 net2947 VPWR VGND sg13g2_buf_8
XFILLER_103_371 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C_sg13g2_nor2_1_Y
+ net3145 net3142 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C
+ VPWR VGND sg13g2_nor2_1
XFILLER_92_704 VPWR VGND sg13g2_decap_4
XFILLER_77_778 VPWR VGND sg13g2_fill_2
XFILLER_65_918 VPWR VGND sg13g2_fill_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_73_940 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.pc_d\[9\]
+ VGND net2304 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xstrb_reg_q\[0\]_sg13g2_nor2_1_A net501 net2730 strb_reg_q\[0\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[293\]_sg13g2_nor3_1_A net1304 net2777 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
XFILLER_72_483 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2829
+ sg13g2_a221oi_1
XFILLER_44_185 VPWR VGND sg13g2_fill_1
XFILLER_33_859 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[16\]_sg13g2_nor2_1_A net546 net2735 shift_reg_q\[16\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] net679 net2617
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2844
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2574 VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ VGND net2582 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_58_4 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[6\]_sg13g2_dfrbpq_1_Q net3197 VGND VPWR net507 shift_reg_q\[6\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2558 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_358 VPWR VGND sg13g2_decap_8
XFILLER_101_308 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0 net3133 i_snitch.i_snitch_regfile.mem\[140\]
+ i_snitch.i_snitch_regfile.mem\[172\] i_snitch.i_snitch_regfile.mem\[204\] i_snitch.i_snitch_regfile.mem\[236\]
+ net3113 i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2632 VPWR i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_67_266 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[75\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2357
+ sg13g2_o21ai_1
XFILLER_49_970 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_X
+ net3095 net2930 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_55_417 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[296\]_sg13g2_o21ai_1_A1 net2937 VPWR i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[296\] net2813 sg13g2_o21ai_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VGND net2588 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_48_491 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1
+ net560 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[435\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net478 net2411 VPWR VGND sg13g2_nand2_1
XFILLER_24_804 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ sg13g2_a21oi_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[224\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[224\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2333 net783 net2903 net2874 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2413
+ sg13g2_o21ai_1
XFILLER_50_155 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2386
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2816 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C net2313 i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.inst_addr_o\[10\] i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D net3250 VGND VPWR data_pvalid_sg13g2_nor2_1_A_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q clknet_leaf_20_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2399
+ sg13g2_o21ai_1
XFILLER_104_168 VPWR VGND sg13g2_decap_8
XFILLER_99_881 VPWR VGND sg13g2_decap_8
XFILLER_59_723 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2597 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_98_391 VPWR VGND sg13g2_decap_8
XFILLER_98_380 VPWR VGND sg13g2_decap_4
XFILLER_58_200 VPWR VGND sg13g2_fill_2
XFILLER_101_875 VPWR VGND sg13g2_decap_8
XFILLER_100_352 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2_sg13g2_nand2b_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2
+ net2516 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2b_1
XFILLER_46_406 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[115\]
+ net2802 sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A net1407 net1410 i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_55_940 VPWR VGND sg13g2_decap_8
Xrebuffer82 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X
+ net114 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C
+ VPWR VGND sg13g2_nand2_1
Xrebuffer71 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ net103 VPWR VGND sg13g2_buf_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1
+ VPWR VGND net3141 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_B1
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xrebuffer60 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X
+ net92 VPWR VGND sg13g2_buf_1
XFILLER_25_20 VPWR VGND sg13g2_fill_1
XFILLER_42_612 VPWR VGND sg13g2_fill_2
Xrebuffer93 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B
+ net125 VPWR VGND sg13g2_buf_2
Xrsp_data_q\[16\]_sg13g2_dfrbpq_1_Q net3234 VGND VPWR rsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[16\] clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_25_42 VPWR VGND sg13g2_fill_2
XFILLER_30_818 VPWR VGND sg13g2_decap_8
XFILLER_42_678 VPWR VGND sg13g2_decap_8
XFILLER_22_391 VPWR VGND sg13g2_fill_1
XFILLER_41_96 VPWR VGND sg13g2_fill_2
Xfanout2700 net2702 net2700 VPWR VGND sg13g2_buf_8
Xfanout2711 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X
+ net2711 VPWR VGND sg13g2_buf_2
XFILLER_2_730 VPWR VGND sg13g2_fill_2
XFILLER_96_328 VPWR VGND sg13g2_decap_4
Xfanout2722 net2726 net2722 VPWR VGND sg13g2_buf_8
Xfanout2744 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y
+ net2744 VPWR VGND sg13g2_buf_8
Xfanout2733 net2734 net2733 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[455\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[244\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net724 net2671 net2875 VPWR VGND sg13g2_a22oi_1
Xfanout2755 net2756 net2755 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2422 sg13g2_a21oi_1
XFILLER_49_200 VPWR VGND sg13g2_decap_4
Xfanout2777 net2778 net2777 VPWR VGND sg13g2_buf_8
Xfanout2788 net2789 net2788 VPWR VGND sg13g2_buf_8
XFILLER_2_796 VPWR VGND sg13g2_decap_8
XFILLER_1_295 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net600 i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2401 net2408 i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_dfrbpq_1_Q_D net2474
+ sg13g2_a221oi_1
Xfanout2766 net2770 net2766 VPWR VGND sg13g2_buf_1
XFILLER_49_255 VPWR VGND sg13g2_decap_4
XFILLER_2_46 VPWR VGND sg13g2_decap_8
Xfanout2799 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_X
+ net2799 VPWR VGND sg13g2_buf_8
XFILLER_92_534 VPWR VGND sg13g2_decap_4
XFILLER_92_545 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[350\] net2951 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[417\]_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_a221oi_1_A1_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_18_675 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2328
+ sg13g2_o21ai_1
XFILLER_60_453 VPWR VGND sg13g2_fill_1
Xheichips25_snitch_wrapper_31 VPWR VGND uio_oe[1] sg13g2_tiehi
XFILLER_21_829 VPWR VGND sg13g2_decap_8
XFILLER_60_475 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q
+ net3244 VGND VPWR net778 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_12_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1_X net2963 VPWR VGND sg13g2_a22oi_1
XFILLER_99_133 VPWR VGND sg13g2_decap_8
XFILLER_82_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_fill_1
XFILLER_101_105 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[349\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[349\] VGND sg13g2_inv_1
XFILLER_96_873 VPWR VGND sg13g2_decap_8
XFILLER_68_564 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ net2705 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ sg13g2_a221oi_1
XFILLER_83_556 VPWR VGND sg13g2_fill_2
XFILLER_71_707 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q_D
+ i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A
+ clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_55_258 VPWR VGND sg13g2_decap_4
XFILLER_102_14 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2570 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_71_718 VPWR VGND sg13g2_fill_2
XFILLER_64_770 VPWR VGND sg13g2_decap_4
XFILLER_52_910 VPWR VGND sg13g2_fill_2
XFILLER_62_29 VPWR VGND sg13g2_fill_1
XFILLER_23_144 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2582 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[475\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_a22oi_1_B2_Y
+ net2325 net634 net2644 net2893 VPWR VGND sg13g2_a22oi_1
XFILLER_106_934 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y net2829 i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2348
+ sg13g2_o21ai_1
XFILLER_79_818 VPWR VGND sg13g2_decap_4
XFILLER_105_499 VPWR VGND sg13g2_fill_2
XFILLER_101_683 VPWR VGND sg13g2_fill_2
XFILLER_101_672 VPWR VGND sg13g2_fill_1
XFILLER_98_1025 VPWR VGND sg13g2_decap_4
XFILLER_87_895 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_fill_1
XFILLER_4_1018 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[147\]
+ i_snitch.i_snitch_regfile.mem\[179\] i_snitch.i_snitch_regfile.mem\[211\] i_snitch.i_snitch_regfile.mem\[243\]
+ net3098 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xdata_pdata\[17\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net730 data_pdata\[17\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y net2717
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_14_144 VPWR VGND sg13g2_fill_2
XFILLER_14_155 VPWR VGND sg13g2_decap_8
XFILLER_42_442 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VGND sg13g2_inv_1
XFILLER_70_784 VPWR VGND sg13g2_fill_1
XFILLER_52_51 VPWR VGND sg13g2_fill_1
XFILLER_14_188 VPWR VGND sg13g2_fill_1
XFILLER_7_822 VPWR VGND sg13g2_decap_8
XFILLER_7_855 VPWR VGND sg13g2_decap_4
XFILLER_7_899 VPWR VGND sg13g2_fill_1
XFILLER_6_387 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B
+ net2636 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xfanout3231 net3232 net3231 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[165\]_sg13g2_nor3_1_A net1239 net2772 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xfanout3220 net3225 net3220 VPWR VGND sg13g2_buf_8
Xfanout3242 net3243 net3242 VPWR VGND sg13g2_buf_8
Xfanout3253 net3259 net3253 VPWR VGND sg13g2_buf_8
Xfanout3264 net3272 net3264 VPWR VGND sg13g2_buf_8
XFILLER_97_659 VPWR VGND sg13g2_decap_8
Xfanout2552 net2553 net2552 VPWR VGND sg13g2_buf_8
Xfanout2541 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y
+ net2541 VPWR VGND sg13g2_buf_8
Xfanout2563 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y
+ net2563 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y net3088
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_2_582 VPWR VGND sg13g2_decap_8
Xfanout3286 net3287 net3286 VPWR VGND sg13g2_buf_8
Xfanout2530 net2534 net2530 VPWR VGND sg13g2_buf_8
Xfanout3275 net3276 net3275 VPWR VGND sg13g2_buf_8
Xfanout3297 net3299 net3297 VPWR VGND sg13g2_buf_8
Xfanout2596 net2597 net2596 VPWR VGND sg13g2_buf_2
Xfanout2574 net2575 net2574 VPWR VGND sg13g2_buf_8
Xfanout2585 net2588 net2585 VPWR VGND sg13g2_buf_2
XFILLER_93_832 VPWR VGND sg13g2_decap_8
XFILLER_77_394 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0 net3013 i_snitch.i_snitch_regfile.mem\[266\]
+ i_snitch.i_snitch_regfile.mem\[298\] i_snitch.i_snitch_regfile.mem\[330\] i_snitch.i_snitch_regfile.mem\[362\]
+ net2986 i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_65_589 VPWR VGND sg13g2_decap_8
XFILLER_52_217 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[495\] clknet_leaf_81_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net1067 net2434 net2247 VPWR VGND sg13g2_a22oi_1
XFILLER_21_604 VPWR VGND sg13g2_fill_2
XFILLER_61_795 VPWR VGND sg13g2_decap_8
XFILLER_61_784 VPWR VGND sg13g2_fill_1
XFILLER_60_261 VPWR VGND sg13g2_decap_4
XFILLER_60_250 VPWR VGND sg13g2_decap_4
XFILLER_33_486 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[86\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[86\]
+ i_snitch.i_snitch_regfile.mem\[118\] net3136 i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2
+ VPWR VGND sg13g2_nor2_1
XFILLER_88_648 VPWR VGND sg13g2_decap_8
XFILLER_84_821 VPWR VGND sg13g2_fill_1
XFILLER_68_361 VPWR VGND sg13g2_decap_8
XFILLER_95_191 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q net3208 VGND VPWR i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[314\] clknet_leaf_117_clk sg13g2_dfrbpq_1
XFILLER_84_898 VPWR VGND sg13g2_decap_8
XFILLER_56_567 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C i_snitch.inst_addr_o\[27\]
+ net106 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_43_228 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2448 net2285 net2409 net1295 VPWR VGND sg13g2_a22oi_1
XFILLER_25_932 VPWR VGND sg13g2_fill_1
XFILLER_36_280 VPWR VGND sg13g2_decap_4
XFILLER_37_792 VPWR VGND sg13g2_decap_4
XFILLER_52_762 VPWR VGND sg13g2_fill_2
XFILLER_19_1026 VPWR VGND sg13g2_fill_2
XFILLER_24_431 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net2695 i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A2
+ net2540 sg13g2_a21oi_1
XFILLER_52_795 VPWR VGND sg13g2_fill_1
XFILLER_106_1018 VPWR VGND sg13g2_decap_8
XFILLER_8_608 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_nand2_1_A_Y net3026 net2998 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_98_14 VPWR VGND sg13g2_decap_8
Xdata_pdata\[13\]_sg13g2_mux2_1_A1 rsp_data_q\[13\] net725 net3049 data_pdata\[13\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_106_720 VPWR VGND sg13g2_decap_8
XFILLER_105_252 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2420 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_65_1024 VPWR VGND sg13g2_decap_4
XFILLER_26_1019 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_A1
+ net1346 VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[438\] net3020 VPWR VGND sg13g2_nand2_1
XFILLER_19_214 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_90_813 VPWR VGND sg13g2_decap_8
XFILLER_74_375 VPWR VGND sg13g2_fill_1
XFILLER_16_943 VPWR VGND sg13g2_decap_8
XFILLER_90_868 VPWR VGND sg13g2_decap_8
XFILLER_62_559 VPWR VGND sg13g2_fill_1
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_72_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[335\] VGND sg13g2_inv_1
XFILLER_15_475 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2757 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
XFILLER_30_445 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1
+ net3083 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[439\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2383 net757 net2647 net2863 VPWR VGND sg13g2_a22oi_1
Xhold608 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net640 sg13g2_dlygate4sd3_1
Xhold619 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\] VPWR
+ VGND net651 sg13g2_dlygate4sd3_1
XFILLER_98_913 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net950 net1069 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[334\] clknet_leaf_78_clk sg13g2_dfrbpq_1
Xfanout3061 net3062 net3061 VPWR VGND sg13g2_buf_8
Xfanout3072 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1_X
+ net3072 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q
+ net3235 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xfanout3050 net3051 net3050 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2448 net2253 net2409 net1234 VPWR VGND sg13g2_a22oi_1
Xfanout3083 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_X
+ net3083 VPWR VGND sg13g2_buf_8
Xfanout2371 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2371 VPWR VGND sg13g2_buf_8
Xfanout3094 net3097 net3094 VPWR VGND sg13g2_buf_8
Xfanout2360 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2360 VPWR VGND sg13g2_buf_8
XFILLER_97_489 VPWR VGND sg13g2_fill_2
Xhold1319 i_snitch.i_snitch_regfile.mem\[299\] VPWR VGND net1351 sg13g2_dlygate4sd3_1
Xfanout2393 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2393 VPWR VGND sg13g2_buf_8
Xfanout2382 net2383 net2382 VPWR VGND sg13g2_buf_8
Xhold1308 i_snitch.i_snitch_regfile.mem\[37\] VPWR VGND net1340 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[43\]_sg13g2_o21ai_1_A1 net3021 VPWR i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[43\] net2994 sg13g2_o21ai_1
XFILLER_93_673 VPWR VGND sg13g2_decap_8
XFILLER_65_353 VPWR VGND sg13g2_fill_1
XFILLER_26_729 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_53_526 VPWR VGND sg13g2_fill_1
XFILLER_19_792 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2557 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_81_879 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[22\]_sg13g2_a22oi_1_A1 shift_reg_q\[22\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[22\] VPWR VGND sg13g2_a22oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B
+ net87 net2928 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_nand3_1
XFILLER_33_250 VPWR VGND sg13g2_fill_1
XFILLER_22_979 VPWR VGND sg13g2_fill_1
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y
+ i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1
+ net3 net645 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]
+ net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_103_701 VPWR VGND sg13g2_decap_8
XFILLER_89_902 VPWR VGND sg13g2_decap_8
XFILLER_88_434 VPWR VGND sg13g2_fill_1
XFILLER_68_28 VPWR VGND sg13g2_fill_2
XFILLER_1_839 VPWR VGND sg13g2_decap_8
XFILLER_103_767 VPWR VGND sg13g2_fill_2
XFILLER_89_979 VPWR VGND sg13g2_decap_8
XFILLER_88_456 VPWR VGND sg13g2_fill_2
XFILLER_102_266 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2696 net37 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ net2541 sg13g2_a21oi_1
Xi_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C
+ i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND sg13g2_nor3_1
XFILLER_84_27 VPWR VGND sg13g2_decap_8
XFILLER_29_545 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y
+ net2610 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B VPWR
+ VGND sg13g2_nor2_1
XFILLER_29_556 VPWR VGND sg13g2_fill_1
XFILLER_71_334 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ net2539 sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_mux2_1_A1
+ net747 net643 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A_sg13g2_nand2b_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A
+ net3093 net40 VPWR VGND sg13g2_nand2b_1
XFILLER_71_345 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[459\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2373 net892 net2679 net2741 VPWR VGND sg13g2_a22oi_1
XFILLER_13_902 VPWR VGND sg13g2_fill_1
XFILLER_13_913 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[354\] clknet_leaf_109_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2352 net1142 net2678 net2890 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_or2_1_X
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net3071 i_snitch.sb_q\[1\] sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2816 i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_X
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 VPWR VGND sg13g2_nor2_1
XFILLER_106_572 VPWR VGND sg13g2_decap_8
XFILLER_79_423 VPWR VGND sg13g2_decap_8
Xrsp_state_d_sg13g2_and2_1_X net4 net3064 rsp_state_d VPWR VGND sg13g2_and2_1
XFILLER_95_938 VPWR VGND sg13g2_decap_8
XFILLER_59_180 VPWR VGND sg13g2_fill_1
XFILLER_12_8 VPWR VGND sg13g2_decap_8
XFILLER_63_813 VPWR VGND sg13g2_decap_8
XFILLER_75_684 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]
+ net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_16_751 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[14\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[14\]
+ i_snitch.inst_addr_o\[14\] clknet_leaf_55_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2866
+ net2898 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y
+ net2923 net2926 net3033 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A
+ VPWR VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ sg13g2_nand4_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N_sg13g2_a21o_1_X
+ net2535 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_req_arb.data_i\[38\] i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N
+ VPWR VGND sg13g2_a21o_1
XFILLER_8_983 VPWR VGND sg13g2_decap_8
XFILLER_7_460 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2641 i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
Xhold427 strb_reg_q\[3\] VPWR VGND net459 sg13g2_dlygate4sd3_1
Xhold416 cnt_q\[2\] VPWR VGND net448 sg13g2_dlygate4sd3_1
Xhold405 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net437 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2 i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_B1 VPWR
+ i_snitch.pc_d\[14\]_sg13g2_o21ai_1_A2_Y VGND i_snitch.inst_addr_o\[14\] i_snitch.pc_d\[14\]
+ sg13g2_o21ai_1
Xhold449 shift_reg_q\[17\] VPWR VGND net481 sg13g2_dlygate4sd3_1
Xhold438 i_snitch.i_snitch_regfile.mem\[321\] VPWR VGND net470 sg13g2_dlygate4sd3_1
XFILLER_86_916 VPWR VGND sg13g2_decap_8
XFILLER_58_607 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_85_404 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2376 net789 net2645 net2740 VPWR VGND sg13g2_a22oi_1
Xhold1105 i_snitch.i_snitch_regfile.mem\[232\] VPWR VGND net1137 sg13g2_dlygate4sd3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q
+ net3240 VGND VPWR net1140 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
Xhold1138 rsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1170
+ sg13g2_dlygate4sd3_1
Xhold1149 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\] VPWR
+ VGND net1181 sg13g2_dlygate4sd3_1
Xhold1116 data_pdata\[8\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net1148 sg13g2_dlygate4sd3_1
Xhold1127 i_snitch.i_snitch_regfile.mem\[467\] VPWR VGND net1159 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net3078 net2537 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ i_snitch.inst_addr_o\[10\] sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[493\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_364 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ net2613 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 VPWR VGND sg13g2_a21o_2
XFILLER_65_183 VPWR VGND sg13g2_fill_2
XFILLER_65_172 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[374\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_0_1010 VPWR VGND sg13g2_decap_8
XFILLER_26_515 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_21_264 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[432\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[70\] VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2501 net2420 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ VGND net2596 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[509\] clknet_leaf_96_clk sg13g2_dfrbpq_1
Xhold972 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold950 i_snitch.i_snitch_regfile.mem\[118\] VPWR VGND net982 sg13g2_dlygate4sd3_1
Xhold961 i_snitch.i_snitch_regfile.mem\[250\] VPWR VGND net993 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y
+ net2618 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_103_542 VPWR VGND sg13g2_fill_2
XFILLER_103_520 VPWR VGND sg13g2_fill_1
XFILLER_89_765 VPWR VGND sg13g2_decap_4
Xhold983 i_snitch.i_snitch_regfile.mem\[108\] VPWR VGND net1015 sg13g2_dlygate4sd3_1
XFILLER_1_636 VPWR VGND sg13g2_decap_8
Xhold994 target_sel_q VPWR VGND net1026 sg13g2_dlygate4sd3_1
XFILLER_103_564 VPWR VGND sg13g2_decap_8
XFILLER_88_253 VPWR VGND sg13g2_fill_2
XFILLER_77_949 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C i_req_arb.data_i\[44\] net2301
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
XFILLER_48_106 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]
+ net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_76_459 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y
+ net44 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ net2509 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2446 VPWR VGND sg13g2_nand2_1
Xi_req_register.data_o\[44\]_sg13g2_o21ai_1_Y i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.data_o\[44\] VGND net3169 i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[102\]
+ net2997 i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_84_470 VPWR VGND sg13g2_decap_4
XFILLER_56_161 VPWR VGND sg13g2_fill_1
XFILLER_44_323 VPWR VGND sg13g2_decap_4
XFILLER_17_537 VPWR VGND sg13g2_fill_1
XFILLER_72_698 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2437 VPWR VGND sg13g2_nand2_1
XFILLER_100_91 VPWR VGND sg13g2_decap_8
XFILLER_9_747 VPWR VGND sg13g2_fill_1
XFILLER_8_213 VPWR VGND sg13g2_fill_2
XFILLER_12_286 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[499\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2271 net2367 net1325 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2892 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2
+ net2507 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_5_942 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2542 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q net3274 VGND VPWR i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[394\] clknet_leaf_101_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y
+ net96 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1
+ VPWR VGND sg13g2_nor3_1
XFILLER_79_264 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[183\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net1078 net2648 net2775 VPWR VGND sg13g2_a22oi_1
XFILLER_67_437 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_82_418 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_and2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_and2_1
XFILLER_78_1001 VPWR VGND sg13g2_decap_8
XFILLER_63_621 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B_sg13g2_nor2_1_Y
+ net2592 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_90_440 VPWR VGND sg13g2_fill_1
XFILLER_35_356 VPWR VGND sg13g2_fill_2
XFILLER_91_996 VPWR VGND sg13g2_decap_8
XFILLER_90_473 VPWR VGND sg13g2_fill_2
XFILLER_23_529 VPWR VGND sg13g2_fill_1
XFILLER_44_890 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1
+ net772 net586 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
XFILLER_102_1010 VPWR VGND sg13g2_decap_8
XFILLER_79_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2432 net2245 net2319 net1161 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[451\] VGND sg13g2_inv_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]
+ net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[213\] clknet_leaf_98_clk sg13g2_dfrbpq_1
XFILLER_105_14 VPWR VGND sg13g2_decap_8
XFILLER_85_201 VPWR VGND sg13g2_fill_2
XFILLER_100_534 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net3180 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]
+ sg13g2_o21ai_1
XFILLER_85_212 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2434 VPWR VGND sg13g2_nand2_1
XFILLER_100_567 VPWR VGND sg13g2_fill_1
XFILLER_67_971 VPWR VGND sg13g2_decap_4
XFILLER_82_930 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2710 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xstrb_reg_q\[2\]_sg13g2_a21oi_1_A1 VGND VPWR net517 net3043 strb_reg_q\[2\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[2\]_sg13g2_a21oi_1_A1_B1 sg13g2_a21oi_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2
+ VPWR VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_Y
+ net2759 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[288\]_sg13g2_dfrbpq_1_Q_D VGND net2315 net2522
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[250\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2957
+ i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2962
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y net49 net2312 net2751 i_snitch.pc_d\[0\]_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_6_706 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1_A1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_B2
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2862
+ net2694 VPWR VGND sg13g2_nand2_1
Xrebuffer387 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1 net419 VPWR VGND sg13g2_buf_1
XFILLER_30_54 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net123 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X net2496 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_2_901 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[336\]_sg13g2_nand2_1_A_1 i_snitch.i_snitch_regfile.mem\[336\]_sg13g2_nand2_1_A_1_Y
+ i_snitch.i_snitch_regfile.mem\[336\] net2951 VPWR VGND sg13g2_nand2_1
XFILLER_104_851 VPWR VGND sg13g2_decap_8
Xfanout2915 net2917 net2915 VPWR VGND sg13g2_buf_8
Xfanout2926 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y
+ net2926 VPWR VGND sg13g2_buf_8
Xfanout2937 net2938 net2937 VPWR VGND sg13g2_buf_8
Xhold780 i_snitch.i_snitch_regfile.mem\[63\] VPWR VGND net812 sg13g2_dlygate4sd3_1
Xfanout2904 data_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y net2904 VPWR
+ VGND sg13g2_buf_8
Xhold791 i_snitch.i_snitch_regfile.mem\[200\] VPWR VGND net823 sg13g2_dlygate4sd3_1
XFILLER_103_350 VPWR VGND sg13g2_decap_8
Xfanout2959 net2960 net2959 VPWR VGND sg13g2_buf_8
XFILLER_49_415 VPWR VGND sg13g2_decap_8
XFILLER_2_978 VPWR VGND sg13g2_decap_8
Xfanout2948 net2949 net2948 VPWR VGND sg13g2_buf_8
XFILLER_89_595 VPWR VGND sg13g2_fill_2
XFILLER_49_426 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[83\]_sg13g2_mux2_1_A0_X net3100 net2824 i_snitch.i_snitch_regfile.mem\[51\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net978 net2454 net2271 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_Y net2979 net2842 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_92_738 VPWR VGND sg13g2_fill_2
XFILLER_64_429 VPWR VGND sg13g2_fill_2
XFILLER_45_621 VPWR VGND sg13g2_fill_2
XFILLER_18_824 VPWR VGND sg13g2_fill_1
XFILLER_29_161 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_a22oi_1_B2_Y
+ net2405 net672 net2473 net2272 VPWR VGND sg13g2_a22oi_1
XFILLER_33_838 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ net88 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2_1_Y
+ net2564 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N
+ VPWR VGND sg13g2_nor2_1
XFILLER_72_495 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]
+ net3170 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_41_871 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2580 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_71_61 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[233\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[233\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_9_544 VPWR VGND sg13g2_fill_1
XFILLER_13_573 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1223 net2492 net1200 VPWR VGND sg13g2_a22oi_1
XFILLER_99_304 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B
+ VGND VPWR i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y sg13g2_nor4_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2705 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_inv_1_A
+ net768 i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_A2 VPWR VGND sg13g2_inv_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ net2612 VPWR VGND sg13g2_a22oi_1
XFILLER_96_91 VPWR VGND sg13g2_decap_4
XFILLER_64_952 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2347
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ net2610 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2843
+ sg13g2_a221oi_1
XFILLER_36_687 VPWR VGND sg13g2_fill_1
XFILLER_90_270 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2475 i_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2436 net2874 i_snitch.i_snitch_regfile.mem\[228\]_sg13g2_dfrbpq_1_Q_D net2907
+ sg13g2_a221oi_1
XFILLER_35_175 VPWR VGND sg13g2_fill_1
XFILLER_52_1026 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2498 net2418 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A
+ VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2461
+ net2513 net2901 net2741 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net987 net2451 net2285 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2483 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[363\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2392
+ sg13g2_o21ai_1
XFILLER_104_147 VPWR VGND sg13g2_decap_8
XFILLER_99_860 VPWR VGND sg13g2_decap_8
XFILLER_59_713 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[358\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net1102 net2899 net2881 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] net662 net2617
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_101_854 VPWR VGND sg13g2_decap_8
XFILLER_100_331 VPWR VGND sg13g2_decap_8
XFILLER_58_267 VPWR VGND sg13g2_decap_4
XFILLER_47_919 VPWR VGND sg13g2_fill_1
XFILLER_74_727 VPWR VGND sg13g2_decap_8
XFILLER_73_215 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[72\]
+ net2842 i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q net3271 VGND VPWR i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[253\] clknet_leaf_92_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1 net3091 VPWR i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[420\] net2811 sg13g2_o21ai_1
Xrebuffer61 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2
+ net93 VPWR VGND sg13g2_buf_1
Xrebuffer72 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ net104 VPWR VGND sg13g2_buf_1
Xrebuffer50 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ net82 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
Xrebuffer83 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ net115 VPWR VGND sg13g2_buf_1
XFILLER_81_292 VPWR VGND sg13g2_fill_1
XFILLER_14_326 VPWR VGND sg13g2_decap_4
XFILLER_27_698 VPWR VGND sg13g2_fill_1
XFILLER_30_808 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_Y
+ VGND net67 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ sg13g2_o21ai_1
Xclkbuf_leaf_115_clk clknet_5_5__leaf_clk clknet_leaf_115_clk VPWR VGND sg13g2_buf_8
XFILLER_41_189 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y
+ net3176 net563 VPWR VGND sg13g2_nand2b_1
XFILLER_6_503 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2_sg13g2_nand3_1_C
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2
+ net2569 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2968 i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
Xfanout2701 net2702 net2701 VPWR VGND sg13g2_buf_1
Xfanout2712 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X
+ net2712 VPWR VGND sg13g2_buf_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_96_307 VPWR VGND sg13g2_decap_8
Xfanout2745 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y
+ net2745 VPWR VGND sg13g2_buf_8
Xfanout2723 net2726 net2723 VPWR VGND sg13g2_buf_1
Xfanout2734 net2737 net2734 VPWR VGND sg13g2_buf_8
XFILLER_2_775 VPWR VGND sg13g2_decap_8
XFILLER_104_692 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
Xfanout2756 net2763 net2756 VPWR VGND sg13g2_buf_2
Xdata_pdata\[0\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B net3153 data_pdata\[0\]_sg13g2_mux2_1_A0_X
+ data_pdata\[0\]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_1_263 VPWR VGND sg13g2_fill_1
XFILLER_2_25 VPWR VGND sg13g2_decap_8
Xfanout2767 net2770 net2767 VPWR VGND sg13g2_buf_8
Xfanout2778 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X
+ net2778 VPWR VGND sg13g2_buf_8
Xfanout2789 net2790 net2789 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2608 net2570 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ net2561 sg13g2_a21oi_1
Xi_snitch.pc_d\[20\]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y_sg13g2_and2_1_A i_snitch.pc_d\[20\]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[23\]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1_Y i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B
+ net3084 net2536 VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1
+ net596 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_80_719 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]_sg13g2_dfrbpq_1_Q
+ net3199 VGND VPWR net611 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[91\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[91\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net1038 net2451 net2253 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net690 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2402 net2485 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D net2474
+ sg13g2_a221oi_1
XFILLER_33_679 VPWR VGND sg13g2_fill_1
Xheichips25_snitch_wrapper_32 VPWR VGND uio_oe[0] sg13g2_tiehi
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y
+ net2758 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2 VPWR VGND sg13g2_nand2_1
XFILLER_60_498 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_106_clk clknet_5_24__leaf_clk clknet_leaf_106_clk VPWR VGND sg13g2_buf_8
XFILLER_20_307 VPWR VGND sg13g2_fill_2
XFILLER_32_189 VPWR VGND sg13g2_fill_2
XFILLER_70_4 VPWR VGND sg13g2_decap_4
XFILLER_9_385 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net1021 net2469 net2255 VPWR VGND sg13g2_a22oi_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2_sg13g2_nand2_1_Y i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2
+ i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_112 VPWR VGND sg13g2_decap_8
XFILLER_88_808 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[273\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_102_607 VPWR VGND sg13g2_decap_4
XFILLER_99_178 VPWR VGND sg13g2_decap_8
XFILLER_96_852 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_29_919 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[379\]
+ net3116 i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_nor2b_1_B_N_Y
+ sg13g2_a21oi_1
XFILLER_28_407 VPWR VGND sg13g2_decap_8
XFILLER_95_395 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2b_1_Y
+ net40 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2b_1
XFILLER_51_410 VPWR VGND sg13g2_fill_2
XFILLER_12_808 VPWR VGND sg13g2_decap_8
XFILLER_24_668 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[408\] clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_51_487 VPWR VGND sg13g2_decap_4
XFILLER_11_329 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_20_885 VPWR VGND sg13g2_fill_2
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
XFILLER_106_913 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2592 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_105_478 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B_Y
+ net645 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_59_510 VPWR VGND sg13g2_decap_8
XFILLER_101_640 VPWR VGND sg13g2_fill_1
XFILLER_87_874 VPWR VGND sg13g2_decap_8
XFILLER_59_554 VPWR VGND sg13g2_fill_2
XFILLER_59_543 VPWR VGND sg13g2_decap_8
Xcnt_q\[2\]_sg13g2_dfrbpq_1_Q net3184 VGND VPWR net450 cnt_q\[2\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
XFILLER_101_662 VPWR VGND sg13g2_fill_1
XFILLER_98_1004 VPWR VGND sg13g2_decap_8
XFILLER_59_576 VPWR VGND sg13g2_decap_8
XFILLER_46_215 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2414
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A_X
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B_X
+ VPWR VGND sg13g2_and4_1
Xstrb_reg_q\[0\]_sg13g2_a22oi_1_A1_B1_sg13g2_nor2_1_Y i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y
+ req_data_valid_sg13g2_o21ai_1_Y_B1 strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B1 VPWR VGND
+ sg13g2_nor2_1
XFILLER_74_579 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[76\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[76\] net2991 VPWR VGND sg13g2_nand2_1
XFILLER_46_259 VPWR VGND sg13g2_fill_2
XFILLER_27_451 VPWR VGND sg13g2_decap_8
XFILLER_54_281 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_fill_2
XFILLER_15_635 VPWR VGND sg13g2_decap_4
XFILLER_27_495 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2390 net1130 net2687 net3041 VPWR VGND sg13g2_a22oi_1
XFILLER_11_852 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q net3222 VGND VPWR i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[293\] clknet_leaf_111_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nand3_1
Xfanout3210 net3211 net3210 VPWR VGND sg13g2_buf_8
Xfanout3221 net3222 net3221 VPWR VGND sg13g2_buf_8
Xfanout3243 net3248 net3243 VPWR VGND sg13g2_buf_8
Xfanout3232 net3249 net3232 VPWR VGND sg13g2_buf_8
Xfanout2520 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X
+ net2520 VPWR VGND sg13g2_buf_8
Xfanout3254 net3258 net3254 VPWR VGND sg13g2_buf_8
Xfanout3265 net3272 net3265 VPWR VGND sg13g2_buf_8
Xfanout2542 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X
+ net2542 VPWR VGND sg13g2_buf_8
Xfanout2553 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C_Y
+ net2553 VPWR VGND sg13g2_buf_8
Xfanout2531 net2534 net2531 VPWR VGND sg13g2_buf_1
Xfanout3287 net3301 net3287 VPWR VGND sg13g2_buf_8
Xfanout3276 net3282 net3276 VPWR VGND sg13g2_buf_8
Xfanout3298 net3299 net3298 VPWR VGND sg13g2_buf_8
Xfanout2575 net2576 net2575 VPWR VGND sg13g2_buf_2
Xfanout2586 net2587 net2586 VPWR VGND sg13g2_buf_8
Xfanout2564 net2568 net2564 VPWR VGND sg13g2_buf_8
XFILLER_78_863 VPWR VGND sg13g2_decap_4
Xfanout2597 net2598 net2597 VPWR VGND sg13g2_buf_1
XFILLER_93_822 VPWR VGND sg13g2_fill_1
XFILLER_93_800 VPWR VGND sg13g2_decap_8
XFILLER_78_896 VPWR VGND sg13g2_decap_8
XFILLER_65_535 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q net3309 VGND VPWR i_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[428\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_93_888 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_Y
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2b_1
XFILLER_46_771 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[217\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net857 net2439 net2266 VPWR VGND sg13g2_a22oi_1
XFILLER_18_462 VPWR VGND sg13g2_fill_1
XFILLER_93_92 VPWR VGND sg13g2_decap_8
XFILLER_52_229 VPWR VGND sg13g2_decap_8
XFILLER_34_933 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q net3289 VGND VPWR i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[112\] clknet_leaf_89_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1 VPWR VGND net3103 net2823
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[32\]
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y net2826 sg13g2_a221oi_1
XFILLER_20_148 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0 net3137 i_snitch.i_snitch_regfile.mem\[151\]
+ i_snitch.i_snitch_regfile.mem\[183\] i_snitch.i_snitch_regfile.mem\[215\] i_snitch.i_snitch_regfile.mem\[247\]
+ net3111 i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_nand2_1_A_Y net3099 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
Xshift_reg_q\[11\]_sg13g2_dfrbpq_1_Q net3195 VGND VPWR net520 shift_reg_q\[11\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2600 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_103_949 VPWR VGND sg13g2_decap_8
XFILLER_102_448 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[108\]
+ net2808 sg13g2_o21ai_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ net2550 VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ VGND net2747 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
XFILLER_68_395 VPWR VGND sg13g2_fill_2
XFILLER_28_215 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[161\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net464 net2342 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[321\]_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_B1
+ i_snitch.i_snitch_regfile.mem\[321\]_sg13g2_o21ai_1_A1_Y VGND sg13g2_inv_1
XFILLER_84_877 VPWR VGND sg13g2_decap_8
XFILLER_83_387 VPWR VGND sg13g2_decap_8
XFILLER_71_549 VPWR VGND sg13g2_fill_2
XFILLER_24_454 VPWR VGND sg13g2_fill_1
XFILLER_25_966 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2
+ VPWR VGND net2699 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1
+ net2544 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_605 VPWR VGND sg13g2_fill_1
XFILLER_51_284 VPWR VGND sg13g2_fill_2
XFILLER_40_947 VPWR VGND sg13g2_fill_1
XFILLER_7_108 VPWR VGND sg13g2_decap_8
XFILLER_22_22 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A net1407 i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_20_671 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_fill_1
XFILLER_106_743 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.i_snitch_regfile.mem\[448\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[448\] clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_3_314 VPWR VGND sg13g2_fill_2
XFILLER_105_231 VPWR VGND sg13g2_decap_8
XFILLER_3_369 VPWR VGND sg13g2_fill_1
XFILLER_106_787 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[237\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net1144 net2690 net2876 VPWR VGND sg13g2_a22oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B
+ VPWR VGND i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
XFILLER_102_982 VPWR VGND sg13g2_decap_8
XFILLER_75_822 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[90\]
+ i_snitch.i_snitch_regfile.mem\[122\] net3119 i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1 net3017 i_snitch.i_snitch_regfile.mem\[141\]
+ i_snitch.i_snitch_regfile.mem\[173\] i_snitch.i_snitch_regfile.mem\[205\] i_snitch.i_snitch_regfile.mem\[237\]
+ net2988 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_101_492 VPWR VGND sg13g2_fill_2
XFILLER_93_129 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[280\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[280\] net3029 VPWR VGND sg13g2_nand2_1
XFILLER_47_41 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[132\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_90_803 VPWR VGND sg13g2_fill_2
XFILLER_75_899 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_and2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1 VPWR VGND net3099 net2821
+ i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[34\]
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y net2824 sg13g2_a221oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2549 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B
+ net2556 sg13g2_a21oi_1
XFILLER_90_847 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\] net2622 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_16_911 VPWR VGND sg13g2_decap_4
XFILLER_27_270 VPWR VGND sg13g2_fill_1
XFILLER_103_91 VPWR VGND sg13g2_decap_8
XFILLER_27_292 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[11\] net873 net2914 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net537 net2493 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2
+ net2551 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[323\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[323\] net2948 VPWR VGND sg13g2_nand2_1
XFILLER_31_969 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ net2486 i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_7_675 VPWR VGND sg13g2_fill_1
Xhold609 i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y VPWR VGND net641 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2558 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xfanout3040 net3042 net3040 VPWR VGND sg13g2_buf_8
Xfanout3073 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X
+ net3073 VPWR VGND sg13g2_buf_8
Xfanout3062 rsp_state_q_sg13g2_nor2_1_A_Y net3062 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[312\] VGND sg13g2_inv_1
Xfanout3051 net3052 net3051 VPWR VGND sg13g2_buf_8
XFILLER_3_892 VPWR VGND sg13g2_decap_8
XFILLER_98_969 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[29\]_sg13g2_dfrbpq_1_Q net3240 VGND VPWR rsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[29\] clknet_leaf_39_clk sg13g2_dfrbpq_2
Xfanout3084 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_X
+ net3084 VPWR VGND sg13g2_buf_1
Xfanout2361 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2361 VPWR VGND sg13g2_buf_8
Xfanout3095 net3097 net3095 VPWR VGND sg13g2_buf_2
Xfanout2350 net2351 net2350 VPWR VGND sg13g2_buf_8
Xfanout2372 net2376 net2372 VPWR VGND sg13g2_buf_8
Xfanout2394 net2398 net2394 VPWR VGND sg13g2_buf_8
Xhold1309 i_snitch.i_snitch_regfile.mem\[386\] VPWR VGND net1341 sg13g2_dlygate4sd3_1
Xfanout2383 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2383 VPWR VGND sg13g2_buf_8
XFILLER_38_502 VPWR VGND sg13g2_decap_8
XFILLER_38_513 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[404\] net3029 VPWR VGND sg13g2_nand2_1
XFILLER_53_505 VPWR VGND sg13g2_decap_8
XFILLER_81_858 VPWR VGND sg13g2_decap_8
XFILLER_80_313 VPWR VGND sg13g2_decap_8
XFILLER_19_782 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VGND net2704 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[468\] clknet_leaf_61_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[442\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[442\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net510 net2384 VPWR VGND sg13g2_nand2_1
XFILLER_21_446 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1_sg13g2_and4_1_X
+ net3035 net2925 net2922 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1
+ VPWR VGND sg13g2_and4_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1 net3021 i_snitch.i_snitch_regfile.mem\[143\]
+ i_snitch.i_snitch_regfile.mem\[175\] i_snitch.i_snitch_regfile.mem\[207\] i_snitch.i_snitch_regfile.mem\[239\]
+ net2992 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[152\] clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_1_818 VPWR VGND sg13g2_decap_8
XFILLER_89_958 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y
+ VGND net2717 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_102_245 VPWR VGND sg13g2_decap_8
XFILLER_88_446 VPWR VGND sg13g2_decap_4
XFILLER_84_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_95_clk clknet_5_17__leaf_clk clknet_leaf_95_clk VPWR VGND sg13g2_buf_8
XFILLER_71_324 VPWR VGND sg13g2_fill_1
XFILLER_16_229 VPWR VGND sg13g2_decap_4
XFILLER_52_571 VPWR VGND sg13g2_fill_1
XFILLER_25_785 VPWR VGND sg13g2_decap_8
XFILLER_40_711 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q
+ net3237 VGND VPWR net646 i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B
+ clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_40_799 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0 net3126 i_snitch.i_snitch_regfile.mem\[158\]
+ i_snitch.i_snitch_regfile.mem\[190\] i_snitch.i_snitch_regfile.mem\[222\] i_snitch.i_snitch_regfile.mem\[254\]
+ net3106 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_95_917 VPWR VGND sg13g2_decap_8
XFILLER_88_980 VPWR VGND sg13g2_decap_8
XFILLER_0_884 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X
+ VPWR VGND sg13g2_and4_1
Xclkbuf_leaf_86_clk clknet_5_22__leaf_clk clknet_leaf_86_clk VPWR VGND sg13g2_buf_8
XFILLER_47_332 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q net3280 VGND VPWR i_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[488\] clknet_leaf_74_clk sg13g2_dfrbpq_1
XFILLER_90_666 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_a22oi_1_B2_Y
+ net2323 net691 net2433 net2269 VPWR VGND sg13g2_a22oi_1
XFILLER_43_571 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2604 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1 net3021 i_snitch.i_snitch_regfile.mem\[145\]
+ i_snitch.i_snitch_regfile.mem\[177\] i_snitch.i_snitch_regfile.mem\[209\] i_snitch.i_snitch_regfile.mem\[241\]
+ net2994 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_15_295 VPWR VGND sg13g2_fill_1
XFILLER_31_722 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q net3317 VGND VPWR i_snitch.i_snitch_regfile.mem\[172\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[172\] clknet_leaf_68_clk sg13g2_dfrbpq_1
XFILLER_30_243 VPWR VGND sg13g2_decap_8
XFILLER_8_940 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_10_clk clknet_5_3__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold406 i_snitch.i_snitch_regfile.mem\[432\] VPWR VGND net438 sg13g2_dlygate4sd3_1
Xhold417 cnt_q\[2\]_sg13g2_a21oi_1_B1_Y VPWR VGND net449 sg13g2_dlygate4sd3_1
XFILLER_99_91 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1 net3009 i_snitch.i_snitch_regfile.mem\[393\]
+ i_snitch.i_snitch_regfile.mem\[425\] i_snitch.i_snitch_regfile.mem\[457\] i_snitch.i_snitch_regfile.mem\[489\]
+ net2982 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xhold428 strb_reg_q\[3\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net460 sg13g2_dlygate4sd3_1
Xhold439 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\] VPWR
+ VGND net471 sg13g2_dlygate4sd3_1
XFILLER_98_722 VPWR VGND sg13g2_decap_4
XFILLER_98_755 VPWR VGND sg13g2_fill_2
XFILLER_98_744 VPWR VGND sg13g2_decap_8
Xhold1106 i_snitch.i_snitch_regfile.mem\[300\] VPWR VGND net1138 sg13g2_dlygate4sd3_1
XFILLER_78_490 VPWR VGND sg13g2_decap_4
Xhold1117 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\] VPWR
+ VGND net1149 sg13g2_dlygate4sd3_1
Xhold1128 i_snitch.i_snitch_lsu.metadata_q\[4\] VPWR VGND net1160 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q net3209 VGND VPWR i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[307\] clknet_leaf_117_clk sg13g2_dfrbpq_1
Xhold1139 i_snitch.i_snitch_regfile.mem\[316\] VPWR VGND net1171 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_77_clk clknet_5_22__leaf_clk clknet_leaf_77_clk VPWR VGND sg13g2_buf_8
XFILLER_65_140 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2920
+ sg13g2_a221oi_1
XFILLER_38_354 VPWR VGND sg13g2_fill_1
XFILLER_94_994 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_Y i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
XFILLER_39_899 VPWR VGND sg13g2_fill_2
XFILLER_55_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2728 shift_reg_q\[25\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[21\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[21\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_34_571 VPWR VGND sg13g2_decap_4
XFILLER_62_891 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[67\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nor3_1_A_Y net2451 net2782 i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_dfrbpq_1_Q_D
+ net2909 sg13g2_a221oi_1
XFILLER_79_17 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2499 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_102_7 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2715 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0 net3134 i_snitch.i_snitch_regfile.mem\[396\]
+ i_snitch.i_snitch_regfile.mem\[428\] i_snitch.i_snitch_regfile.mem\[460\] i_snitch.i_snitch_regfile.mem\[492\]
+ net3113 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold940 i_snitch.i_snitch_regfile.mem\[222\] VPWR VGND net972 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A
+ VPWR VGND sg13g2_xor2_1
Xhold973 i_snitch.i_snitch_regfile.mem\[247\] VPWR VGND net1005 sg13g2_dlygate4sd3_1
Xhold962 i_snitch.i_snitch_regfile.mem\[84\] VPWR VGND net994 sg13g2_dlygate4sd3_1
XFILLER_1_615 VPWR VGND sg13g2_decap_8
Xhold951 i_snitch.i_snitch_regfile.mem\[464\] VPWR VGND net983 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[297\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2685 net2778 net2320 net1280 VPWR VGND sg13g2_a22oi_1
Xhold984 i_snitch.i_snitch_regfile.mem\[221\] VPWR VGND net1016 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold995 target_sel_q_sg13g2_dfrbpq_1_Q_D VPWR VGND net1027 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y
+ sg13g2_a21oi_2
XFILLER_62_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_608 VPWR VGND sg13g2_decap_4
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_95_49 VPWR VGND sg13g2_decap_8
XFILLER_76_438 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1 net2999 i_snitch.i_snitch_regfile.mem\[147\]
+ i_snitch.i_snitch_regfile.mem\[179\] i_snitch.i_snitch_regfile.mem\[211\] i_snitch.i_snitch_regfile.mem\[243\]
+ net2973 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net60 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2_Y
+ net2564 sg13g2_a21oi_1
Xclkbuf_leaf_68_clk clknet_5_27__leaf_clk clknet_leaf_68_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[192\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[192\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_85_983 VPWR VGND sg13g2_decap_8
XFILLER_17_505 VPWR VGND sg13g2_fill_1
XFILLER_72_677 VPWR VGND sg13g2_decap_8
Xdata_pdata\[24\]_sg13g2_mux2_1_A1 rsp_data_q\[24\] net927 net3051 data_pdata\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_44_379 VPWR VGND sg13g2_fill_2
XFILLER_32_519 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[40\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_12_232 VPWR VGND sg13g2_decap_4
XFILLER_12_254 VPWR VGND sg13g2_decap_8
XFILLER_100_70 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[376\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[344\]_sg13g2_inv_1_A_Y net3137 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net485 net2373 VPWR VGND sg13g2_nand2_1
XFILLER_5_921 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[327\] clknet_leaf_117_clk sg13g2_dfrbpq_1
XFILLER_5_998 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_106_392 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[116\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[116\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net1060 net2671 net2871 VPWR VGND sg13g2_a22oi_1
XFILLER_69_72 VPWR VGND sg13g2_decap_4
XFILLER_69_61 VPWR VGND sg13g2_fill_2
Xi_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1
+ net2487 i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_68_928 VPWR VGND sg13g2_decap_8
XFILLER_68_917 VPWR VGND sg13g2_fill_1
XFILLER_67_416 VPWR VGND sg13g2_decap_4
XFILLER_95_736 VPWR VGND sg13g2_decap_4
XFILLER_0_681 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_59_clk clknet_5_31__leaf_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
XFILLER_48_663 VPWR VGND sg13g2_fill_1
XFILLER_76_983 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1
+ net3179 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] VPWR
+ VGND sg13g2_nand2_1
XFILLER_36_869 VPWR VGND sg13g2_decap_4
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[15\]_sg13g2_a22oi_1_A1 shift_reg_q\[15\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_mux2_1_A1_1_X
+ net3055 net3045 net461 VPWR VGND sg13g2_a22oi_1
XFILLER_91_975 VPWR VGND sg13g2_decap_8
XFILLER_90_452 VPWR VGND sg13g2_decap_8
XFILLER_23_508 VPWR VGND sg13g2_fill_1
XFILLER_90_496 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q
+ net3231 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_43_390 VPWR VGND sg13g2_fill_2
XFILLER_31_552 VPWR VGND sg13g2_decap_8
XFILLER_105_819 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1 net3005 i_snitch.i_snitch_regfile.mem\[149\]
+ i_snitch.i_snitch_regfile.mem\[181\] i_snitch.i_snitch_regfile.mem\[213\] i_snitch.i_snitch_regfile.mem\[245\]
+ net2978 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_104_329 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_A2
+ net2542 VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2
+ net41 i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ sg13g2_a21oi_1
XFILLER_85_224 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[88\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_nand2b_1_A_N_Y
+ net3030 i_snitch.i_snitch_regfile.mem\[88\] VPWR VGND sg13g2_nand2b_1
XFILLER_22_1001 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1 net3017 i_snitch.i_snitch_regfile.mem\[397\]
+ i_snitch.i_snitch_regfile.mem\[429\] i_snitch.i_snitch_regfile.mem\[461\] i_snitch.i_snitch_regfile.mem\[493\]
+ net2988 i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[60\] clknet_leaf_101_clk sg13g2_dfrbpq_1
XFILLER_39_685 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2422 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_53_121 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
XFILLER_82_986 VPWR VGND sg13g2_decap_8
XFILLER_54_688 VPWR VGND sg13g2_fill_1
XFILLER_42_828 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[347\] clknet_leaf_117_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2423 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1_sg13g2_inv_1_Y i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1
+ net1119 VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[136\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2352 net752 net2643 net2887 VPWR VGND sg13g2_a22oi_1
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_104_830 VPWR VGND sg13g2_decap_8
Xfanout2916 net2917 net2916 VPWR VGND sg13g2_buf_1
Xfanout2927 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net2927 VPWR VGND sg13g2_buf_8
Xhold781 i_snitch.i_snitch_regfile.mem\[351\] VPWR VGND net813 sg13g2_dlygate4sd3_1
Xhold770 i_snitch.i_snitch_regfile.mem\[383\] VPWR VGND net802 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_1_423 VPWR VGND sg13g2_fill_1
Xfanout2905 data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2905 VPWR VGND
+ sg13g2_buf_8
Xfanout2949 net111 net2949 VPWR VGND sg13g2_buf_8
Xfanout2938 net2939 net2938 VPWR VGND sg13g2_buf_8
XFILLER_1_467 VPWR VGND sg13g2_fill_2
Xhold792 data_pdata\[10\] VPWR VGND net824 sg13g2_dlygate4sd3_1
XFILLER_89_585 VPWR VGND sg13g2_fill_1
XFILLER_65_909 VPWR VGND sg13g2_fill_1
XFILLER_58_972 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ net2571 VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VGND i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_44_121 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2440 VPWR VGND sg13g2_nand2_1
XFILLER_45_677 VPWR VGND sg13g2_fill_2
Xdata_pdata\[1\]_sg13g2_dfrbpq_1_Q net3196 VGND VPWR net735 data_pdata\[1\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1
+ net2489 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C
+ VPWR VGND sg13g2_and3_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[424\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2379
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[309\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2778
+ net2670 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1 net3020 i_snitch.i_snitch_regfile.mem\[399\]
+ i_snitch.i_snitch_regfile.mem\[431\] i_snitch.i_snitch_regfile.mem\[463\] i_snitch.i_snitch_regfile.mem\[495\]
+ net2992 i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2845
+ sg13g2_a221oi_1
XFILLER_4_283 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[80\] clknet_leaf_88_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_96_70 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_83_706 VPWR VGND sg13g2_fill_1
XFILLER_67_235 VPWR VGND sg13g2_decap_4
XFILLER_95_577 VPWR VGND sg13g2_fill_1
XFILLER_67_268 VPWR VGND sg13g2_fill_1
XFILLER_55_419 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[367\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net937 net2447 net2246 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y_sg13g2_inv_1_A
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_inv_2
XFILLER_91_761 VPWR VGND sg13g2_decap_8
XFILLER_63_441 VPWR VGND sg13g2_decap_8
XFILLER_51_603 VPWR VGND sg13g2_fill_1
XFILLER_35_132 VPWR VGND sg13g2_decap_4
XFILLER_91_1010 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y
+ VPWR VGND sg13g2_nor4_1
XFILLER_91_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2357
+ sg13g2_o21ai_1
XFILLER_51_658 VPWR VGND sg13g2_decap_8
XFILLER_23_349 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1
+ net573 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_nand2_1_A_Y net3031 net2997 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_104_126 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0
+ VGND net2607 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_101_833 VPWR VGND sg13g2_decap_8
XFILLER_100_310 VPWR VGND sg13g2_decap_8
XFILLER_86_511 VPWR VGND sg13g2_fill_1
XFILLER_86_500 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_A1
+ net1372 VGND sg13g2_inv_1
XFILLER_74_706 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[27\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[27\]
+ i_snitch.inst_addr_o\[27\] clknet_leaf_52_clk sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ net2969 VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B
+ VGND i_snitch.sb_q\[10\] i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
XFILLER_100_387 VPWR VGND sg13g2_fill_1
XFILLER_86_588 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ sg13g2_o21ai_1
XFILLER_92_28 VPWR VGND sg13g2_decap_8
Xrebuffer51 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ net83 VPWR VGND sg13g2_buf_1
Xrebuffer62 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y
+ net94 VPWR VGND sg13g2_buf_1
Xrebuffer73 net3183 net105 VPWR VGND sg13g2_buf_1
Xrebuffer40 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ net72 VPWR VGND sg13g2_buf_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1153 net2495 net1291 VPWR VGND sg13g2_a22oi_1
XFILLER_54_463 VPWR VGND sg13g2_fill_1
XFILLER_54_441 VPWR VGND sg13g2_fill_2
Xrebuffer84 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X
+ net116 VPWR VGND sg13g2_buf_1
XFILLER_25_44 VPWR VGND sg13g2_fill_1
XFILLER_26_187 VPWR VGND sg13g2_decap_8
XFILLER_42_614 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ net2716 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_23_850 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X net2509
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_10_533 VPWR VGND sg13g2_fill_1
XFILLER_22_382 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nand3_1_Y
+ net2926 net2925 net2922 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nand3_1
XFILLER_41_98 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[387\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[387\] clknet_leaf_112_clk sg13g2_dfrbpq_1
Xfanout2702 net2703 net2702 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[379\]
+ net2800 i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xfanout2713 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X
+ net2713 VPWR VGND sg13g2_buf_1
Xfanout2724 net2726 net2724 VPWR VGND sg13g2_buf_8
Xfanout2735 net2736 net2735 VPWR VGND sg13g2_buf_2
XFILLER_2_754 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[176\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2444 net2263 net2344 net1275 VPWR VGND sg13g2_a22oi_1
XFILLER_104_682 VPWR VGND sg13g2_fill_2
Xfanout2746 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y
+ net2746 VPWR VGND sg13g2_buf_1
XFILLER_89_371 VPWR VGND sg13g2_decap_8
XFILLER_77_511 VPWR VGND sg13g2_fill_2
Xfanout2757 net2758 net2757 VPWR VGND sg13g2_buf_8
XFILLER_49_224 VPWR VGND sg13g2_fill_1
Xfanout2779 net2781 net2779 VPWR VGND sg13g2_buf_8
Xfanout2768 net2770 net2768 VPWR VGND sg13g2_buf_8
XFILLER_1_297 VPWR VGND sg13g2_fill_1
XFILLER_38_909 VPWR VGND sg13g2_fill_1
XFILLER_106_91 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2706 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_92_503 VPWR VGND sg13g2_fill_1
XFILLER_46_942 VPWR VGND sg13g2_fill_2
XFILLER_46_931 VPWR VGND sg13g2_decap_8
XFILLER_18_622 VPWR VGND sg13g2_decap_8
XFILLER_18_633 VPWR VGND sg13g2_fill_2
XFILLER_92_569 VPWR VGND sg13g2_fill_2
XFILLER_45_441 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y
+ net2581 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_75_1027 VPWR VGND sg13g2_fill_2
XFILLER_60_422 VPWR VGND sg13g2_decap_4
XFILLER_60_400 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y net2309
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B
+ net93 VPWR VGND sg13g2_nand2_1
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_9_364 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ VGND net2573 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q net3289 VGND VPWR i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[206\] clknet_leaf_88_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X_sg13g2_a21o_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_B
+ VPWR VGND sg13g2_a21o_1
XFILLER_96_831 VPWR VGND sg13g2_decap_8
XFILLER_95_330 VPWR VGND sg13g2_fill_1
XFILLER_83_525 VPWR VGND sg13g2_decap_8
XFILLER_55_238 VPWR VGND sg13g2_decap_4
XFILLER_102_49 VPWR VGND sg13g2_decap_8
XFILLER_91_580 VPWR VGND sg13g2_decap_4
XFILLER_64_794 VPWR VGND sg13g2_fill_1
XFILLER_63_271 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.sb_q\[1\] net2826 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ net2823 sg13g2_a21oi_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A
+ net39 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor4_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_A i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B
+ i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[502\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net1109 net2651 net2857 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[4\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C net3153 data_pdata\[12\]_sg13g2_nor2b_1_A_Y
+ data_pdata\[4\]_sg13g2_nor2_1_B_Y data_pdata\[4\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_106_969 VPWR VGND sg13g2_decap_8
XFILLER_105_413 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2552 VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[76\]_sg13g2_mux2_1_A0_X net3113 net2829 i_snitch.i_snitch_regfile.mem\[44\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2779
+ net2694 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[44\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net1082 net2692 net2769 VPWR VGND sg13g2_a22oi_1
XFILLER_59_500 VPWR VGND sg13g2_fill_1
XFILLER_87_853 VPWR VGND sg13g2_decap_8
XFILLER_59_533 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[303\] VGND sg13g2_inv_1
XFILLER_101_685 VPWR VGND sg13g2_fill_1
XFILLER_100_140 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[503\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[503\]
+ net3137 i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
XFILLER_100_184 VPWR VGND sg13g2_decap_8
XFILLER_86_385 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2348
+ sg13g2_o21ai_1
XFILLER_74_547 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ net2566 sg13g2_a21oi_1
XFILLER_43_945 VPWR VGND sg13g2_fill_2
XFILLER_14_124 VPWR VGND sg13g2_fill_1
XFILLER_15_658 VPWR VGND sg13g2_decap_8
XFILLER_15_669 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[226\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_42_433 VPWR VGND sg13g2_decap_8
XFILLER_70_775 VPWR VGND sg13g2_decap_8
XFILLER_43_989 VPWR VGND sg13g2_fill_2
XFILLER_35_1000 VPWR VGND sg13g2_fill_2
XFILLER_42_488 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_mux2_1_A1
+ net1069 net552 net2237 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.sb_q\[3\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[3\] i_snitch.sb_q\[3\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2738
+ net2897 VPWR VGND sg13g2_nand2_1
XFILLER_30_639 VPWR VGND sg13g2_fill_2
XFILLER_10_352 VPWR VGND sg13g2_decap_4
XFILLER_6_301 VPWR VGND sg13g2_decap_4
XFILLER_7_846 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A
+ net2549 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ net72 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_6_356 VPWR VGND sg13g2_decap_4
Xfanout3200 net3205 net3200 VPWR VGND sg13g2_buf_8
Xfanout3211 net3226 net3211 VPWR VGND sg13g2_buf_8
Xfanout3222 net3224 net3222 VPWR VGND sg13g2_buf_8
XFILLER_97_617 VPWR VGND sg13g2_decap_8
Xfanout3244 net3247 net3244 VPWR VGND sg13g2_buf_8
Xfanout2510 net2511 net2510 VPWR VGND sg13g2_buf_8
Xfanout3233 net3236 net3233 VPWR VGND sg13g2_buf_8
Xfanout3255 net3258 net3255 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ state sg13g2_a21oi_1
XFILLER_105_980 VPWR VGND sg13g2_decap_8
Xfanout2554 net2556 net2554 VPWR VGND sg13g2_buf_8
Xfanout2543 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X
+ net2543 VPWR VGND sg13g2_buf_8
Xfanout2532 net2534 net2532 VPWR VGND sg13g2_buf_8
Xfanout2521 i_snitch.consec_pc\[0\]_sg13g2_a22oi_1_A1_Y net2521 VPWR VGND sg13g2_buf_8
Xfanout3266 net3272 net3266 VPWR VGND sg13g2_buf_8
Xfanout3288 net3301 net3288 VPWR VGND sg13g2_buf_8
Xfanout3277 net3281 net3277 VPWR VGND sg13g2_buf_8
XFILLER_35_8 VPWR VGND sg13g2_decap_8
Xfanout3299 net3300 net3299 VPWR VGND sg13g2_buf_8
Xfanout2587 net2588 net2587 VPWR VGND sg13g2_buf_8
Xfanout2565 net2567 net2565 VPWR VGND sg13g2_buf_8
Xfanout2576 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y
+ net2576 VPWR VGND sg13g2_buf_8
Xuio_out_sg13g2_inv_1_Y_1 VPWR net11 uio_out_sg13g2_inv_1_Y_1_A VGND sg13g2_inv_1
Xfanout2598 net2599 net2598 VPWR VGND sg13g2_buf_1
XFILLER_77_374 VPWR VGND sg13g2_fill_1
Xcnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A
+ cnt_q\[2\]_sg13g2_nand3_1_A_Y state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 VPWR
+ VGND sg13g2_nor2_1
XFILLER_93_867 VPWR VGND sg13g2_decap_8
XFILLER_92_366 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_37_249 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A
+ VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_80_528 VPWR VGND sg13g2_decap_8
XFILLER_73_580 VPWR VGND sg13g2_fill_2
XFILLER_45_271 VPWR VGND sg13g2_decap_8
XFILLER_33_400 VPWR VGND sg13g2_decap_8
XFILLER_33_411 VPWR VGND sg13g2_fill_1
XFILLER_61_753 VPWR VGND sg13g2_fill_2
XFILLER_61_742 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B
+ net2931 i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_21_606 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand4_1_Y
+ net2925 net2922 net3035 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2354 net765 net2904 net2785 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
XFILLER_9_194 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2883
+ net2650 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net523 net2355 VPWR VGND sg13g2_nand2_1
XFILLER_88_617 VPWR VGND sg13g2_decap_8
XFILLER_103_928 VPWR VGND sg13g2_decap_8
XFILLER_84_801 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q net3320 VGND VPWR i_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[246\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_3_91 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[413\]_sg13g2_o21ai_1_A1 net3094 VPWR i_snitch.i_snitch_regfile.mem\[413\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[413\] net2814 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2458 VPWR VGND sg13g2_nand2_1
XFILLER_84_856 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2490 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_o21ai_1
XFILLER_56_525 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1 net2999 i_snitch.i_snitch_regfile.mem\[411\]
+ i_snitch.i_snitch_regfile.mem\[443\] i_snitch.i_snitch_regfile.mem\[475\] i_snitch.i_snitch_regfile.mem\[507\]
+ net2973 i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_926 VPWR VGND sg13g2_decap_4
XFILLER_12_639 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_105_210 VPWR VGND sg13g2_decap_8
XFILLER_98_49 VPWR VGND sg13g2_decap_8
XFILLER_106_766 VPWR VGND sg13g2_decap_8
XFILLER_105_287 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ sg13g2_o21ai_1
XFILLER_102_961 VPWR VGND sg13g2_decap_8
XFILLER_59_363 VPWR VGND sg13g2_decap_4
XFILLER_101_471 VPWR VGND sg13g2_decap_4
XFILLER_74_311 VPWR VGND sg13g2_fill_1
XFILLER_59_396 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[84\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2356 net994 net2672 net2787 VPWR VGND sg13g2_a22oi_1
XFILLER_103_70 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_xnor2_1
XFILLER_72_1019 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.inst_addr_o\[30\] net2721 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_C1 sg13g2_a21oi_1
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_Y
+ VGND net2718 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_43_797 VPWR VGND sg13g2_fill_2
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_31_948 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[266\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[266\] clknet_leaf_101_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
Xfanout3030 net3031 net3030 VPWR VGND sg13g2_buf_8
XFILLER_98_948 VPWR VGND sg13g2_decap_8
Xfanout3063 net3064 net3063 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q
+ net3238 VGND VPWR net874 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_1
Xfanout3052 target_sel_q_sg13g2_nand2_1_B_Y net3052 VPWR VGND sg13g2_buf_8
XFILLER_3_871 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y net2956
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xfanout3041 net3042 net3041 VPWR VGND sg13g2_buf_8
Xfanout3085 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1_X
+ net3085 VPWR VGND sg13g2_buf_8
Xfanout3074 net3075 net3074 VPWR VGND sg13g2_buf_8
Xfanout2340 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2340 VPWR VGND sg13g2_buf_8
Xfanout3096 net3097 net3096 VPWR VGND sg13g2_buf_8
Xfanout2351 net2352 net2351 VPWR VGND sg13g2_buf_8
Xfanout2362 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2362 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y
+ VPWR VGND sg13g2_nor3_1
Xfanout2373 net2375 net2373 VPWR VGND sg13g2_buf_8
Xfanout2395 net2397 net2395 VPWR VGND sg13g2_buf_8
Xfanout2384 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2384 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[26\] net758 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_77_182 VPWR VGND sg13g2_decap_4
XFILLER_93_653 VPWR VGND sg13g2_fill_2
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
XFILLER_65_377 VPWR VGND sg13g2_decap_8
XFILLER_34_720 VPWR VGND sg13g2_decap_8
XFILLER_80_336 VPWR VGND sg13g2_decap_4
Xtarget_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A target_sel_q_sg13g2_nand2b_1_A_N_Y
+ target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_18_293 VPWR VGND sg13g2_decap_8
XFILLER_22_915 VPWR VGND sg13g2_fill_2
XFILLER_33_241 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VGND net2712 i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ sg13g2_o21ai_1
XFILLER_22_959 VPWR VGND sg13g2_decap_4
XFILLER_33_296 VPWR VGND sg13g2_decap_4
XFILLER_30_992 VPWR VGND sg13g2_fill_1
XFILLER_88_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_o21ai_1_A1_Y net3088 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y sg13g2_a221oi_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2 VPWR
+ VGND net2757 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 net3074 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y
+ net2853 sg13g2_a221oi_1
XFILLER_89_937 VPWR VGND sg13g2_decap_8
XFILLER_88_414 VPWR VGND sg13g2_fill_2
XFILLER_103_769 VPWR VGND sg13g2_fill_1
XFILLER_102_224 VPWR VGND sg13g2_decap_8
XFILLER_88_458 VPWR VGND sg13g2_fill_1
XFILLER_97_992 VPWR VGND sg13g2_decap_8
XFILLER_96_491 VPWR VGND sg13g2_decap_4
XFILLER_84_631 VPWR VGND sg13g2_fill_1
XFILLER_57_823 VPWR VGND sg13g2_fill_2
XFILLER_56_322 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2764
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_57_878 VPWR VGND sg13g2_decap_8
XFILLER_95_1008 VPWR VGND sg13g2_decap_8
XFILLER_84_697 VPWR VGND sg13g2_decap_8
XFILLER_25_731 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ net2637 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ net2725 i_snitch.inst_addr_o\[15\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[358\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C net3163 i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nand2b_1_B_Y
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y VPWR VGND sg13g2_nor3_2
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[286\] clknet_leaf_93_clk sg13g2_dfrbpq_1
XFILLER_40_734 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C_sg13g2_nand4_1_Y
+ net3083 net3077 net3085 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C
+ VPWR VGND net3079 sg13g2_nand4_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q
+ net3243 VGND VPWR net832 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q
+ net3190 VGND VPWR net621 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_32_1025 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.inst_addr_o\[20\]
+ net2525 VPWR VGND sg13g2_xnor2_1
XFILLER_106_530 VPWR VGND sg13g2_decap_8
XFILLER_4_668 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_167 VPWR VGND sg13g2_fill_1
XFILLER_3_189 VPWR VGND sg13g2_fill_2
XFILLER_0_863 VPWR VGND sg13g2_decap_8
XFILLER_58_85 VPWR VGND sg13g2_fill_2
XFILLER_75_675 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y net110 i_snitch.i_snitch_regfile.mem\[264\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[296\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_47_366 VPWR VGND sg13g2_fill_1
XFILLER_35_528 VPWR VGND sg13g2_fill_1
XFILLER_63_859 VPWR VGND sg13g2_fill_2
XFILLER_62_325 VPWR VGND sg13g2_fill_1
XFILLER_16_720 VPWR VGND sg13g2_decap_8
XFILLER_16_731 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[289\]_sg13g2_a221oi_1_A1 VPWR VGND net2920 net3094
+ i_snitch.i_snitch_regfile.mem\[257\] i_snitch.i_snitch_regfile.mem\[289\] i_snitch.i_snitch_regfile.mem\[289\]_sg13g2_a221oi_1_A1_Y
+ net2825 sg13g2_a221oi_1
XFILLER_90_678 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1
+ net44 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[105\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_15_241 VPWR VGND sg13g2_decap_8
XFILLER_95_7 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] net3179 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_12_970 VPWR VGND sg13g2_decap_8
Xhold407 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\] VPWR
+ VGND net439 sg13g2_dlygate4sd3_1
Xhold418 cnt_q\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net450 sg13g2_dlygate4sd3_1
XFILLER_99_70 VPWR VGND sg13g2_decap_8
Xhold429 shift_reg_q\[15\] VPWR VGND net461 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1
+ VGND VPWR net3134 net2849 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ sg13g2_a21oi_1
Xhold1107 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] VPWR
+ VGND net1139 sg13g2_dlygate4sd3_1
XFILLER_85_439 VPWR VGND sg13g2_fill_1
XFILLER_85_428 VPWR VGND sg13g2_decap_8
XFILLER_66_631 VPWR VGND sg13g2_decap_4
Xhold1129 i_snitch.i_snitch_regfile.mem\[318\] VPWR VGND net1161 sg13g2_dlygate4sd3_1
Xhold1118 i_snitch.i_snitch_regfile.mem\[262\] VPWR VGND net1150 sg13g2_dlygate4sd3_1
XFILLER_94_973 VPWR VGND sg13g2_decap_8
XFILLER_39_856 VPWR VGND sg13g2_decap_8
XFILLER_65_196 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_19_580 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[206\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2391 net975 net2663 net3042 VPWR VGND sg13g2_a22oi_1
XFILLER_53_358 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y
+ net3079 net3081 net3085 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y net489 VPWR i_snitch.sb_d\[4\] VGND net2293 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\] net2623 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_21_299 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[308\] VGND sg13g2_inv_1
Xhold930 i_snitch.i_snitch_regfile.mem\[89\] VPWR VGND net962 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ VGND sg13g2_inv_1
XFILLER_88_200 VPWR VGND sg13g2_decap_4
Xhold941 i_snitch.i_snitch_regfile.mem\[480\] VPWR VGND net973 sg13g2_dlygate4sd3_1
Xhold952 i_snitch.i_snitch_regfile.mem\[219\] VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold963 data_pdata\[11\] VPWR VGND net995 sg13g2_dlygate4sd3_1
XFILLER_103_544 VPWR VGND sg13g2_fill_1
Xhold974 i_snitch.i_snitch_regfile.mem\[249\] VPWR VGND net1006 sg13g2_dlygate4sd3_1
XFILLER_0_126 VPWR VGND sg13g2_decap_8
Xhold996 i_snitch.i_snitch_regfile.mem\[234\] VPWR VGND net1028 sg13g2_dlygate4sd3_1
Xhold985 i_snitch.i_snitch_regfile.mem\[493\] VPWR VGND net1017 sg13g2_dlygate4sd3_1
XFILLER_95_28 VPWR VGND sg13g2_decap_8
XFILLER_77_918 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net2543 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[125\] clknet_leaf_101_clk sg13g2_dfrbpq_1
XFILLER_85_962 VPWR VGND sg13g2_decap_8
XFILLER_69_491 VPWR VGND sg13g2_fill_1
XFILLER_72_601 VPWR VGND sg13g2_fill_1
XFILLER_57_675 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_inv_1_A_Y
+ net2622 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_45_815 VPWR VGND sg13g2_fill_2
XFILLER_84_494 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xi_req_arb.data_i\[44\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.pc_d\[9\] i_req_arb.data_i\[44\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
XFILLER_44_369 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[176\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[20\]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1 i_snitch.pc_d\[20\]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[20\]_sg13g2_or2_1_B_X i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2_Y
+ net419 i_snitch.inst_addr_o\[28\] VPWR VGND sg13g2_a22oi_1
Xshift_reg_q\[24\]_sg13g2_dfrbpq_1_Q net3229 VGND VPWR net530 shift_reg_q\[24\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_9_727 VPWR VGND sg13g2_decap_8
XFILLER_13_756 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_B1
+ VGND VPWR net2716 net47 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VGND net2711 i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
XFILLER_8_248 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 net2629 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_977 VPWR VGND sg13g2_decap_8
XFILLER_106_371 VPWR VGND sg13g2_decap_8
XFILLER_95_759 VPWR VGND sg13g2_fill_2
XFILLER_79_288 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[19\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VGND sg13g2_inv_1
XFILLER_0_660 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[334\] net2951 VPWR VGND sg13g2_nand2_1
XFILLER_48_642 VPWR VGND sg13g2_fill_2
XFILLER_75_450 VPWR VGND sg13g2_fill_2
XFILLER_47_152 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0 net3120 i_snitch.i_snitch_regfile.mem\[405\]
+ i_snitch.i_snitch_regfile.mem\[437\] i_snitch.i_snitch_regfile.mem\[469\] i_snitch.i_snitch_regfile.mem\[501\]
+ net3101 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_91_954 VPWR VGND sg13g2_decap_8
XFILLER_63_645 VPWR VGND sg13g2_fill_1
XFILLER_90_475 VPWR VGND sg13g2_fill_1
XFILLER_63_689 VPWR VGND sg13g2_fill_1
XFILLER_63_678 VPWR VGND sg13g2_decap_4
XFILLER_16_550 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2500 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_62_199 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[422\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[422\]
+ net3014 i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_a21oi_1_A1_Y net2986 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q_D VGND net2315 net2242
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[438\] VGND sg13g2_inv_1
XFILLER_85_1018 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[145\] clknet_leaf_81_clk sg13g2_dfrbpq_1
XFILLER_104_308 VPWR VGND sg13g2_decap_8
XFILLER_98_531 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[127\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2837 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_58_406 VPWR VGND sg13g2_fill_1
XFILLER_100_514 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y VGND
+ VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y sg13g2_a21oi_1
XFILLER_105_49 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[453\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[453\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[453\] net2947 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2447 net2886 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_dfrbpq_1_Q_D net2909
+ sg13g2_a221oi_1
XFILLER_82_965 VPWR VGND sg13g2_decap_8
Xdata_pdata\[31\]_sg13g2_a21oi_1_A2 VGND VPWR net3160 data_pdata\[31\] data_pdata\[31\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[23\]_sg13g2_nor2b_1_B_N_Y sg13g2_a21oi_1
XFILLER_26_358 VPWR VGND sg13g2_fill_1
XFILLER_81_497 VPWR VGND sg13g2_fill_2
XFILLER_81_486 VPWR VGND sg13g2_decap_8
XFILLER_41_317 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[441\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[441\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2463 net2266 net2384 net1186 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[251\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xfanout2928 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net2928 VPWR VGND sg13g2_buf_8
Xfanout2917 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y net2917 VPWR
+ VGND sg13g2_buf_8
Xhold782 i_snitch.i_snitch_regfile.mem\[76\] VPWR VGND net814 sg13g2_dlygate4sd3_1
Xhold760 i_snitch.i_snitch_regfile.mem\[433\] VPWR VGND net792 sg13g2_dlygate4sd3_1
XFILLER_2_936 VPWR VGND sg13g2_decap_8
Xfanout2906 data_pdata\[21\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2906 VPWR VGND
+ sg13g2_buf_8
Xhold771 data_pdata\[21\] VPWR VGND net803 sg13g2_dlygate4sd3_1
XFILLER_89_553 VPWR VGND sg13g2_decap_4
XFILLER_77_704 VPWR VGND sg13g2_fill_1
Xfanout2939 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net2939 VPWR VGND sg13g2_buf_8
Xhold793 data_pdata\[10\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net825 sg13g2_dlygate4sd3_1
XFILLER_104_886 VPWR VGND sg13g2_decap_8
XFILLER_103_385 VPWR VGND sg13g2_decap_8
XFILLER_76_214 VPWR VGND sg13g2_decap_8
XFILLER_76_203 VPWR VGND sg13g2_fill_2
XFILLER_7_1018 VPWR VGND sg13g2_decap_8
XFILLER_58_940 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2
+ net41 sg13g2_a21oi_2
XFILLER_57_483 VPWR VGND sg13g2_fill_2
XFILLER_45_645 VPWR VGND sg13g2_fill_2
XFILLER_45_623 VPWR VGND sg13g2_fill_1
XFILLER_73_987 VPWR VGND sg13g2_fill_1
XFILLER_72_453 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[165\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[165\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_513 VPWR VGND sg13g2_decap_4
XFILLER_40_361 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X
+ net55 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_xor2_1
XFILLER_9_579 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1
+ VPWR VGND net2631 net2565 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C
+ net2548 sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B net2429
+ net2516 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2
+ VGND net2745 net2548 sg13g2_o21ai_1
XFILLER_68_715 VPWR VGND sg13g2_decap_4
XFILLER_45_1013 VPWR VGND sg13g2_decap_8
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1
+ net3072 VPWR VGND sg13g2_inv_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_83_729 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2417 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_24_818 VPWR VGND sg13g2_decap_8
XFILLER_24_829 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[461\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net1044 net2689 net2742 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_and3_1
XFILLER_32_851 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2758 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
XFILLER_52_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_361 VPWR VGND sg13g2_decap_8
XFILLER_84_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2347
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2502 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_105_628 VPWR VGND sg13g2_decap_8
XFILLER_104_105 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nor2_1_Y
+ net3083 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C
+ VPWR VGND sg13g2_nor2_1
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_101_812 VPWR VGND sg13g2_decap_8
XFILLER_99_895 VPWR VGND sg13g2_decap_8
XFILLER_58_214 VPWR VGND sg13g2_decap_8
XFILLER_86_556 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.data_o\[44\]_sg13g2_o21ai_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2497 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_A1 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[185\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[185\] clknet_leaf_116_clk sg13g2_dfrbpq_1
XFILLER_101_889 VPWR VGND sg13g2_decap_8
XFILLER_100_366 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2392
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y
+ VGND VPWR net2581 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ net2577 sg13g2_a21oi_1
Xrebuffer30 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1 net62 VPWR VGND sg13g2_buf_1
Xrebuffer41 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_X
+ net73 VPWR VGND sg13g2_buf_1
Xrebuffer63 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y
+ net95 VPWR VGND sg13g2_buf_2
Xrebuffer52 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ net84 VPWR VGND sg13g2_buf_1
Xrebuffer85 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X
+ net117 VPWR VGND sg13g2_buf_1
Xrebuffer74 net2311 net106 VPWR VGND sg13g2_buf_8
XFILLER_14_317 VPWR VGND sg13g2_fill_2
XFILLER_27_689 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q net3276 VGND VPWR i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[33\] clknet_leaf_104_clk sg13g2_dfrbpq_1
XFILLER_10_501 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[303\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_a22oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2264
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1
+ net2751 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_10_567 VPWR VGND sg13g2_decap_8
XFILLER_41_66 VPWR VGND sg13g2_fill_2
XFILLER_6_538 VPWR VGND sg13g2_fill_1
XFILLER_68_1024 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[122\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2836 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[68\]_sg13g2_nand2b_1_A_N_Y
+ net3032 i_snitch.i_snitch_regfile.mem\[68\] VPWR VGND sg13g2_nand2b_1
Xfanout2703 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X
+ net2703 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2411 net1007 net2690 net2870 VPWR VGND sg13g2_a22oi_1
Xhold590 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\] VPWR
+ VGND net622 sg13g2_dlygate4sd3_1
Xfanout2725 net2726 net2725 VPWR VGND sg13g2_buf_8
Xfanout2736 net2737 net2736 VPWR VGND sg13g2_buf_1
Xfanout2714 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2714 VPWR VGND sg13g2_buf_8
Xstrb_reg_q\[3\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net460 strb_reg_q\[3\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
Xfanout2747 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y
+ net2747 VPWR VGND sg13g2_buf_8
XFILLER_89_383 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y
+ net2949 net40 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nor2_1
Xfanout2758 net2763 net2758 VPWR VGND sg13g2_buf_8
Xfanout2769 net2770 net2769 VPWR VGND sg13g2_buf_8
XFILLER_106_70 VPWR VGND sg13g2_decap_8
XFILLER_103_182 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_77_556 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C net2312 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[6\]_sg13g2_o21ai_1_A2_A1 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]
+ net3178 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_66_30 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C
+ net2564 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X
+ VPWR VGND sg13g2_or3_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2590 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_nand2_1
Xhold1290 rsp_data_q\[6\] VPWR VGND net1322 sg13g2_dlygate4sd3_1
XFILLER_75_1006 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2545 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2426 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q
+ net3192 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
XFILLER_61_968 VPWR VGND sg13g2_fill_2
XFILLER_14_851 VPWR VGND sg13g2_fill_2
XFILLER_13_350 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1
+ net544 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xi_req_arb.data_i\[42\]_sg13g2_inv_1_A net1196 i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y
+ VPWR VGND sg13g2_inv_4
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2321
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[193\]
+ i_snitch.i_snitch_regfile.mem\[225\] net3013 i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[372\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[372\] net2806 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q net3303 VGND VPWR i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[511\] clknet_leaf_72_clk sg13g2_dfrbpq_1
XFILLER_99_147 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2691 net2780 net2318 net1138 VPWR VGND sg13g2_a22oi_1
XFILLER_101_119 VPWR VGND sg13g2_decap_8
XFILLER_95_320 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2335
+ sg13g2_o21ai_1
XFILLER_96_887 VPWR VGND sg13g2_decap_8
XFILLER_55_206 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q net3266 VGND VPWR i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[53\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_102_28 VPWR VGND sg13g2_decap_8
XFILLER_52_935 VPWR VGND sg13g2_decap_8
XFILLER_91_592 VPWR VGND sg13g2_decap_4
XFILLER_52_968 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[301\]
+ net3017 i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_a21oi_1_A1_Y net2988 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y
+ net3093 i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_mux2_1_A0_1_X net3107 net2920 i_snitch.i_snitch_regfile.mem\[129\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_32_681 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ VGND i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B_sg13g2_inv_1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B
+ net92 VGND sg13g2_inv_1
XFILLER_11_14 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_o21ai_1_A1 net3017 VPWR i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[49\] net2988 sg13g2_o21ai_1
XFILLER_106_948 VPWR VGND sg13g2_decap_8
XFILLER_99_681 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[307\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2777
+ net2674 VPWR VGND sg13g2_nand2_1
XFILLER_86_331 VPWR VGND sg13g2_fill_2
XFILLER_86_320 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
XFILLER_86_353 VPWR VGND sg13g2_decap_8
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[182\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2341
+ sg13g2_o21ai_1
XFILLER_19_409 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_B1 VPWR
+ i_snitch.sb_d\[11\] VGND net2292 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_27_420 VPWR VGND sg13g2_fill_2
XFILLER_28_932 VPWR VGND sg13g2_decap_8
XFILLER_28_943 VPWR VGND sg13g2_fill_1
XFILLER_42_412 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[11\]_sg13g2_nor2_1_A net519 net2731 shift_reg_q\[11\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_35_1023 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[320\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2402 net717 net2904 net2795 VPWR VGND sg13g2_a22oi_1
XFILLER_10_386 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_C1
+ net2626 sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2481 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[73\] clknet_leaf_50_clk sg13g2_dfrbpq_1
Xfanout3212 net3213 net3212 VPWR VGND sg13g2_buf_8
Xfanout3201 net3202 net3201 VPWR VGND sg13g2_buf_8
Xfanout3245 net3247 net3245 VPWR VGND sg13g2_buf_8
Xfanout3234 net3236 net3234 VPWR VGND sg13g2_buf_8
Xfanout2511 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B_Y
+ net2511 VPWR VGND sg13g2_buf_8
Xfanout2500 net2501 net2500 VPWR VGND sg13g2_buf_8
Xfanout3256 net3258 net3256 VPWR VGND sg13g2_buf_8
Xfanout3223 net3224 net3223 VPWR VGND sg13g2_buf_8
Xfanout2544 net2545 net2544 VPWR VGND sg13g2_buf_8
XFILLER_78_810 VPWR VGND sg13g2_fill_2
Xfanout2533 net2534 net2533 VPWR VGND sg13g2_buf_8
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1 VGND VPWR data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X
+ sg13g2_a21oi_1
Xfanout2522 i_snitch.consec_pc\[0\]_sg13g2_a22oi_1_A1_Y net2522 VPWR VGND sg13g2_buf_8
Xfanout3267 net3268 net3267 VPWR VGND sg13g2_buf_8
Xfanout3289 net3290 net3289 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[262\] VGND sg13g2_inv_1
Xfanout3278 net3281 net3278 VPWR VGND sg13g2_buf_8
Xfanout2555 net2556 net2555 VPWR VGND sg13g2_buf_1
Xfanout2577 net2578 net2577 VPWR VGND sg13g2_buf_8
Xfanout2566 net2567 net2566 VPWR VGND sg13g2_buf_8
Xuio_out_sg13g2_inv_1_Y_2 VPWR net10 uio_out_sg13g2_inv_1_Y_2_A VGND sg13g2_inv_1
Xfanout2588 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ net2588 VPWR VGND sg13g2_buf_1
Xfanout2599 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_X
+ net2599 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2876
+ net2693 VPWR VGND sg13g2_nand2_1
XFILLER_93_846 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2349 net1087 net2447 net2268 VPWR VGND sg13g2_a22oi_1
XFILLER_19_921 VPWR VGND sg13g2_fill_1
XFILLER_92_345 VPWR VGND sg13g2_fill_2
XFILLER_46_751 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_nand4_1_D
+ net3036 net2927 net3147 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ sg13g2_nand4_1
XFILLER_18_497 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[69\]_sg13g2_o21ai_1_A1 net3099 VPWR i_snitch.i_snitch_regfile.mem\[69\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[69\] net3117 sg13g2_o21ai_1
XFILLER_61_776 VPWR VGND sg13g2_fill_1
XFILLER_33_456 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2798
+ net2676 VPWR VGND sg13g2_nand2_1
XFILLER_103_907 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ VGND sg13g2_inv_1
Xi_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y VGND
+ VPWR i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1
+ i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2
+ i_snitch.wake_up_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0 net1122 sg13g2_a21oi_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2707 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]
+ net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ net3076 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_68_342 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_29_729 VPWR VGND sg13g2_fill_2
XFILLER_96_695 VPWR VGND sg13g2_decap_4
XFILLER_84_835 VPWR VGND sg13g2_decap_8
XFILLER_68_397 VPWR VGND sg13g2_fill_1
Xcnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D VGND net500 cnt_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_28_239 VPWR VGND sg13g2_decap_8
XFILLER_83_334 VPWR VGND sg13g2_fill_2
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y
+ VPWR VGND net2924 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1
+ net2744 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_56_559 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[24\]_sg13g2_nor2_1_A net529 net2736 shift_reg_q\[24\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[340\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2403 net864 net2672 net2796 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q net3270 VGND VPWR i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[93\] clknet_leaf_101_clk sg13g2_dfrbpq_1
Xdata_pdata\[0\]_sg13g2_mux2_1_A0 data_pdata\[0\] data_pdata\[8\] net3161 data_pdata\[0\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q
+ net3238 VGND VPWR net992 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
XFILLER_22_35 VPWR VGND sg13g2_fill_2
XFILLER_22_57 VPWR VGND sg13g2_fill_2
XFILLER_106_734 VPWR VGND sg13g2_decap_8
XFILLER_98_28 VPWR VGND sg13g2_decap_8
XFILLER_4_839 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[169\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2343 net1029 net2686 net2773 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2562 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_105_266 VPWR VGND sg13g2_decap_8
XFILLER_102_940 VPWR VGND sg13g2_decap_8
XFILLER_87_640 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[257\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2434
+ net2514 net2902 net2894 VPWR VGND sg13g2_a22oi_1
XFILLER_87_684 VPWR VGND sg13g2_decap_4
XFILLER_19_228 VPWR VGND sg13g2_decap_8
XFILLER_62_529 VPWR VGND sg13g2_fill_2
XFILLER_28_762 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2464 VPWR VGND sg13g2_nand2_1
XFILLER_34_209 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C VPWR VGND sg13g2_or3_1
XFILLER_16_957 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2499 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_242 VPWR VGND sg13g2_decap_8
XFILLER_42_286 VPWR VGND sg13g2_fill_2
XFILLER_11_651 VPWR VGND sg13g2_decap_4
XFILLER_30_459 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q
+ net3227 VGND VPWR net578 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
XFILLER_7_633 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[21\] net833 net2914 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A
+ VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B
+ net3073 sg13g2_o21ai_1
Xfanout3031 net3032 net3031 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR
+ net2531 net2486 i_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D i_snitch.i_snitch_lsu.metadata_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xfanout3020 net3021 net3020 VPWR VGND sg13g2_buf_8
XFILLER_98_927 VPWR VGND sg13g2_decap_8
Xfanout3064 net3067 net3064 VPWR VGND sg13g2_buf_8
XFILLER_3_850 VPWR VGND sg13g2_decap_8
Xfanout3053 net3055 net3053 VPWR VGND sg13g2_buf_8
Xfanout3042 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y net3042 VPWR VGND sg13g2_buf_8
Xfanout3086 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1_1_X
+ net3086 VPWR VGND sg13g2_buf_1
Xfanout3075 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X
+ net3075 VPWR VGND sg13g2_buf_8
Xfanout2341 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2341 VPWR VGND sg13g2_buf_8
Xfanout3097 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_X
+ net3097 VPWR VGND sg13g2_buf_8
Xfanout2330 net2333 net2330 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[360\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2396 net737 net2644 net2882 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y VPWR VGND net2767 sg13g2_nand2b_2
Xfanout2352 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2352 VPWR VGND sg13g2_buf_8
XFILLER_78_673 VPWR VGND sg13g2_fill_1
Xfanout2385 net2386 net2385 VPWR VGND sg13g2_buf_8
Xfanout2396 net2397 net2396 VPWR VGND sg13g2_buf_8
Xfanout2374 net2376 net2374 VPWR VGND sg13g2_buf_8
Xfanout2363 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ net2363 VPWR VGND sg13g2_buf_8
XFILLER_78_684 VPWR VGND sg13g2_fill_1
XFILLER_66_879 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X
+ VPWR VGND sg13g2_xnor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[361\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[361\]
+ net3123 i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_a21oi_1_A1_Y net2946 sg13g2_a21oi_1
XFILLER_21_437 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[189\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2444 net2250 net2344 net1276 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2295 net1384 net2492 net1342 VPWR VGND sg13g2_a22oi_1
XFILLER_103_715 VPWR VGND sg13g2_fill_2
XFILLER_102_203 VPWR VGND sg13g2_decap_8
XFILLER_89_916 VPWR VGND sg13g2_decap_8
XFILLER_103_737 VPWR VGND sg13g2_decap_4
XFILLER_97_971 VPWR VGND sg13g2_decap_8
XFILLER_69_695 VPWR VGND sg13g2_fill_1
XFILLER_29_537 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 net82
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_44_518 VPWR VGND sg13g2_fill_2
XFILLER_37_570 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A_sg13g2_nand2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q
+ net3230 VGND VPWR net640 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[219\] clknet_leaf_119_clk sg13g2_dfrbpq_1
XFILLER_25_743 VPWR VGND sg13g2_decap_4
XFILLER_37_592 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[38\]
+ net2829 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y net2822 sg13g2_a21oi_1
XFILLER_52_562 VPWR VGND sg13g2_decap_8
XFILLER_52_540 VPWR VGND sg13g2_fill_2
XFILLER_80_882 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2764
+ net2674 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1
+ net2586 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[380\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net1173 net2469 net2246 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_647 VPWR VGND sg13g2_decap_8
XFILLER_106_586 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_58_20 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[380\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2884
+ net2656 VPWR VGND sg13g2_nand2_1
XFILLER_0_842 VPWR VGND sg13g2_decap_8
Xcnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B state cnt_q\[2\]_sg13g2_nand3_1_A_Y
+ cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X VPWR VGND sg13g2_and2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]
+ net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_101_280 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1
+ VGND net2604 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_90_613 VPWR VGND sg13g2_decap_4
XFILLER_63_827 VPWR VGND sg13g2_decap_8
XFILLER_28_581 VPWR VGND sg13g2_fill_2
XFILLER_74_96 VPWR VGND sg13g2_fill_1
XFILLER_16_765 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[271\]_sg13g2_o21ai_1_A1 net2937 VPWR i_snitch.i_snitch_regfile.mem\[271\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[271\] net2814 sg13g2_o21ai_1
XFILLER_31_724 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net830 net2454 net2267 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q net3206 VGND VPWR i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[410\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ net2550 VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B
+ VGND net2715 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xdata_pdata\[7\]_sg13g2_mux2_1_A0 data_pdata\[7\] data_pdata\[15\] net3161 data_pdata\[7\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xhold408 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net440 sg13g2_dlygate4sd3_1
XFILLER_8_997 VPWR VGND sg13g2_decap_8
XFILLER_7_474 VPWR VGND sg13g2_decap_4
Xhold419 i_snitch.i_snitch_regfile.mem\[336\] VPWR VGND net451 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
XFILLER_97_256 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[406\]_sg13g2_o21ai_1_A1 net3097 VPWR i_snitch.i_snitch_regfile.mem\[406\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[406\] i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q net3299 VGND VPWR i_snitch.i_snitch_regfile.mem\[239\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[239\] clknet_leaf_81_clk sg13g2_dfrbpq_1
Xtarget_sel_q_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR target_sel_q_sg13g2_nor2_1_A_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_a21oi_1_A2_Y
+ target_sel_q_sg13g2_dfrbpq_1_Q_D target_sel_q_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold1108 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1140 sg13g2_dlygate4sd3_1
XFILLER_85_418 VPWR VGND sg13g2_decap_4
XFILLER_79_993 VPWR VGND sg13g2_decap_8
XFILLER_78_470 VPWR VGND sg13g2_fill_1
Xhold1119 i_snitch.i_snitch_regfile.mem\[153\] VPWR VGND net1151 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[82\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2786
+ net2676 VPWR VGND sg13g2_nand2_1
XFILLER_39_824 VPWR VGND sg13g2_decap_8
XFILLER_39_835 VPWR VGND sg13g2_fill_2
XFILLER_94_952 VPWR VGND sg13g2_decap_8
XFILLER_65_164 VPWR VGND sg13g2_decap_4
XFILLER_54_827 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[237\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_93_495 VPWR VGND sg13g2_decap_8
XFILLER_0_1024 VPWR VGND sg13g2_decap_4
XFILLER_21_212 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_nand2b_1_A_N_Y
+ net118 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\] VPWR
+ VGND sg13g2_nand2b_1
XFILLER_9_80 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2734 shift_reg_q\[26\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[22\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[22\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xshift_reg_q\[1\]_sg13g2_dfrbpq_1_Q net3186 VGND VPWR net536 shift_reg_q\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
Xhold931 i_snitch.i_snitch_regfile.mem\[327\] VPWR VGND net963 sg13g2_dlygate4sd3_1
Xhold920 i_snitch.i_snitch_regfile.mem\[494\] VPWR VGND net952 sg13g2_dlygate4sd3_1
XFILLER_89_713 VPWR VGND sg13g2_fill_2
Xhold953 i_snitch.i_snitch_regfile.mem\[372\] VPWR VGND net985 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[464\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold942 i_snitch.i_snitch_regfile.mem\[174\] VPWR VGND net974 sg13g2_dlygate4sd3_1
Xhold964 data_pdata\[11\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net996 sg13g2_dlygate4sd3_1
Xhold986 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\] VPWR
+ VGND net1018 sg13g2_dlygate4sd3_1
Xhold997 i_snitch.i_snitch_regfile.mem\[169\] VPWR VGND net1029 sg13g2_dlygate4sd3_1
XFILLER_0_105 VPWR VGND sg13g2_decap_8
Xhold975 i_snitch.i_snitch_regfile.mem\[109\] VPWR VGND net1007 sg13g2_dlygate4sd3_1
XFILLER_85_941 VPWR VGND sg13g2_decap_8
XFILLER_57_632 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q net3295 VGND VPWR i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[430\] clknet_leaf_85_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X net1361 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1
+ net2312 i_snitch.pc_d\[6\] VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net1115 net2690 net2786 VPWR VGND sg13g2_a22oi_1
XFILLER_29_356 VPWR VGND sg13g2_fill_2
XFILLER_72_646 VPWR VGND sg13g2_decap_8
XFILLER_72_635 VPWR VGND sg13g2_fill_2
XFILLER_45_849 VPWR VGND sg13g2_decap_8
XFILLER_25_562 VPWR VGND sg13g2_decap_8
XFILLER_40_521 VPWR VGND sg13g2_decap_4
XFILLER_80_690 VPWR VGND sg13g2_fill_2
XFILLER_52_392 VPWR VGND sg13g2_decap_4
XFILLER_60_54 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[267\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[78\]
+ net2844 i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[259\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[259\] clknet_leaf_105_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_5_956 VPWR VGND sg13g2_decap_8
XFILLER_4_411 VPWR VGND sg13g2_fill_1
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_106_350 VPWR VGND sg13g2_decap_8
XFILLER_69_41 VPWR VGND sg13g2_fill_1
XFILLER_4_466 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_A
+ net50 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_67_407 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR VGND sg13g2_a21o_1
XFILLER_78_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a22oi_1_A2 i_snitch.pc_d\[28\]_sg13g2_a22oi_1_A2_Y i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.inst_addr_o\[31\] i_snitch.pc_d\[28\] i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_63_602 VPWR VGND sg13g2_fill_1
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1
+ net2487 i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_91_933 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[11\]_sg13g2_dfrbpq_1_Q net3230 VGND VPWR rsp_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[11\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_47_186 VPWR VGND sg13g2_decap_4
Xi_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B
+ net553 net545 i_snitch.wake_up_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C
+ VPWR VGND sg13g2_and3_1
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_50_307 VPWR VGND sg13g2_fill_2
XFILLER_31_510 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2
+ net2504 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[11\]_sg13g2_a21o_1_A2 i_snitch.pc_d\[11\] i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1
+ i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_B1 i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X VPWR
+ VGND sg13g2_a21o_1
XFILLER_31_598 VPWR VGND sg13g2_decap_4
XFILLER_102_1024 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[450\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[450\] clknet_leaf_110_clk sg13g2_dfrbpq_1
XFILLER_98_510 VPWR VGND sg13g2_fill_1
XFILLER_98_554 VPWR VGND sg13g2_decap_8
XFILLER_105_28 VPWR VGND sg13g2_decap_8
XFILLER_98_576 VPWR VGND sg13g2_decap_8
XFILLER_86_749 VPWR VGND sg13g2_fill_1
XFILLER_39_610 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[415\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[300\] net3024 VPWR VGND sg13g2_nand2_1
XFILLER_82_944 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[279\] clknet_leaf_70_clk sg13g2_dfrbpq_1
XFILLER_35_893 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR net713 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A_Y
+ strb_reg_q\[4\]_sg13g2_a21oi_1_A1_B1 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_2_915 VPWR VGND sg13g2_decap_8
Xhold761 i_snitch.i_snitch_regfile.mem\[399\] VPWR VGND net793 sg13g2_dlygate4sd3_1
Xhold750 i_snitch.i_snitch_regfile.mem\[251\] VPWR VGND net782 sg13g2_dlygate4sd3_1
Xfanout2918 net81 net2918 VPWR VGND sg13g2_buf_8
Xhold772 data_pdata\[21\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net804 sg13g2_dlygate4sd3_1
Xfanout2907 data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2907 VPWR VGND
+ sg13g2_buf_8
XFILLER_104_865 VPWR VGND sg13g2_decap_8
XFILLER_89_565 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[31\]_sg13g2_dfrbpq_1_Q net3239 VGND VPWR rsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[31\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xhold783 i_snitch.i_snitch_regfile.mem\[456\] VPWR VGND net815 sg13g2_dlygate4sd3_1
Xhold794 i_snitch.i_snitch_regfile.mem\[475\] VPWR VGND net826 sg13g2_dlygate4sd3_1
Xfanout2929 net2932 net2929 VPWR VGND sg13g2_buf_8
XFILLER_103_364 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y VPWR
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y
+ VGND i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ net2626 sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C
+ VGND net2837 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_1_469 VPWR VGND sg13g2_fill_1
XFILLER_39_66 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
XFILLER_92_708 VPWR VGND sg13g2_fill_2
XFILLER_29_142 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2759 net2304
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2517 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_73_933 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net41 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_326 VPWR VGND sg13g2_fill_2
XFILLER_44_156 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_118_clk clknet_5_4__leaf_clk clknet_leaf_118_clk VPWR VGND sg13g2_buf_8
Xi_snitch.sb_q\[15\]_sg13g2_dfrbpq_1_Q net3254 VGND VPWR i_snitch.sb_d\[15\] i_snitch.sb_q\[15\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_41_830 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[470\] clknet_leaf_62_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2778
+ i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2605 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_13_598 VPWR VGND sg13g2_fill_2
Xdata_pdata\[13\]_sg13g2_nand2b_1_B data_pdata\[13\]_sg13g2_nand2b_1_B_Y data_pdata\[13\]
+ net3155 VPWR VGND sg13g2_nand2b_1
XFILLER_40_395 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_nor2_1_Y
+ net2922 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B_sg13g2_a21oi_1_A2
+ VGND VPWR net2570 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C
+ net2579 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[425\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2380
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[299\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_48_462 VPWR VGND sg13g2_fill_1
XFILLER_36_602 VPWR VGND sg13g2_fill_1
Xdata_pdata\[12\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR net902 data_pdata\[12\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_48_495 VPWR VGND sg13g2_fill_2
XFILLER_48_484 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VGND net2558 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ sg13g2_o21ai_1
XFILLER_90_240 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2757 net2303
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1 net2517 sg13g2_a221oi_1
Xclkbuf_leaf_109_clk clknet_5_7__leaf_clk clknet_leaf_109_clk VPWR VGND sg13g2_buf_8
XFILLER_90_295 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.inst_addr_o\[22\]
+ net2525 VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0 net3115 i_snitch.i_snitch_regfile.mem\[135\]
+ i_snitch.i_snitch_regfile.mem\[167\] i_snitch.i_snitch_regfile.mem\[199\] i_snitch.i_snitch_regfile.mem\[231\]
+ net3098 i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_32_841 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[168\]_sg13g2_dfrbpq_1_Q_D VGND net2278 net2340
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2530 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2479 VPWR VGND sg13g2_a22oi_1
XFILLER_32_863 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_77_0 VPWR VGND sg13g2_decap_8
XFILLER_105_607 VPWR VGND sg13g2_fill_2
XFILLER_6_70 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[95\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[95\]_sg13g2_nand2b_1_A_N_Y
+ net3027 i_snitch.i_snitch_regfile.mem\[95\] VPWR VGND sg13g2_nand2b_1
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1
+ net555 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
XFILLER_99_874 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2413
+ sg13g2_o21ai_1
XFILLER_98_384 VPWR VGND sg13g2_fill_2
XFILLER_98_373 VPWR VGND sg13g2_decap_8
XFILLER_86_502 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q net3320 VGND VPWR i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[118\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_101_868 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[4\] i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q_D VGND net2281 net2385
+ sg13g2_o21ai_1
XFILLER_100_345 VPWR VGND sg13g2_decap_8
XFILLER_67_771 VPWR VGND sg13g2_fill_1
Xrebuffer20 net51 net52 VPWR VGND sg13g2_buf_1
Xdata_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2714 data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y net3070 sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[490\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[490\] clknet_leaf_102_clk sg13g2_dfrbpq_1
XFILLER_39_484 VPWR VGND sg13g2_fill_2
Xrebuffer42 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[14\]_sg13g2_mux2_1_A1_1_X
+ net74 VPWR VGND sg13g2_buf_1
Xrebuffer64 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_A
+ net96 VPWR VGND sg13g2_buf_2
Xrebuffer53 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A
+ net85 VPWR VGND sg13g2_buf_1
XFILLER_82_763 VPWR VGND sg13g2_fill_2
XFILLER_82_741 VPWR VGND sg13g2_fill_1
Xrebuffer31 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y
+ net63 VPWR VGND sg13g2_buf_1
Xi_req_arb.data_i\[37\]_sg13g2_dfrbpq_1_Q net3253 VGND VPWR i_snitch.pc_d\[2\] i_req_arb.data_i\[37\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_55_988 VPWR VGND sg13g2_decap_8
Xrebuffer86 net3182 net118 VPWR VGND sg13g2_buf_1
Xrebuffer75 net3140 net107 VPWR VGND sg13g2_buf_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B
+ net2744 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B
+ VPWR VGND i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2
+ sg13g2_nand3b_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y
+ VPWR VGND i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_A2 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2496 i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[41\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xshift_reg_q\[17\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net482 shift_reg_q\[17\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR net3096 net2852 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y sg13g2_a21oi_1
XFILLER_22_373 VPWR VGND sg13g2_fill_1
XFILLER_23_896 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_C1 net2637 i_snitch.inst_addr_o\[31\]
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y
+ net2720 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2408 i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2471 net2878 i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q_D net2906
+ sg13g2_a221oi_1
Xrebuffer198 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ net230 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[486\]_sg13g2_o21ai_1_A1 net2964 VPWR i_snitch.i_snitch_regfile.mem\[486\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[486\] net2804 sg13g2_o21ai_1
XFILLER_2_712 VPWR VGND sg13g2_decap_8
XFILLER_104_651 VPWR VGND sg13g2_fill_2
Xfanout2704 net2705 net2704 VPWR VGND sg13g2_buf_8
Xfanout2715 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y
+ net2715 VPWR VGND sg13g2_buf_8
Xfanout2726 net97 net2726 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2421 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[414\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2467 net2244 net2391 net1155 VPWR VGND sg13g2_a22oi_1
Xhold580 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\] VPWR
+ VGND net612 sg13g2_dlygate4sd3_1
Xfanout2748 net2749 net2748 VPWR VGND sg13g2_buf_8
XFILLER_89_362 VPWR VGND sg13g2_fill_2
XFILLER_77_513 VPWR VGND sg13g2_fill_1
Xfanout2759 net2760 net2759 VPWR VGND sg13g2_buf_8
Xhold591 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\] VPWR
+ VGND net623 sg13g2_dlygate4sd3_1
XFILLER_2_789 VPWR VGND sg13g2_fill_2
Xfanout2737 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y net2737
+ VPWR VGND sg13g2_buf_8
XFILLER_103_161 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[12\]_sg13g2_mux2_1_A1 i_snitch.pc_d\[12\]_sg13g2_mux2_1_A1_A0 i_snitch.pc_d\[12\]
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_A1 i_snitch.pc_d\[12\]_sg13g2_mux2_1_A1_X VPWR
+ VGND sg13g2_mux2_1
XFILLER_2_39 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A_Y net2843 i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_92_538 VPWR VGND sg13g2_fill_2
XFILLER_92_527 VPWR VGND sg13g2_decap_8
XFILLER_57_270 VPWR VGND sg13g2_decap_8
Xhold1291 rsp_data_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1323 sg13g2_dlygate4sd3_1
Xhold1280 i_snitch.i_snitch_regfile.mem\[197\] VPWR VGND net1312 sg13g2_dlygate4sd3_1
XFILLER_18_679 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2365
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ net2560 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_mux2_1
XFILLER_13_384 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ VGND i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_2
XFILLER_12_1002 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[305\]_sg13g2_o21ai_1_A1 net2937 VPWR i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[305\] net2812 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[345\] net2948 VPWR VGND sg13g2_nand2_1
XFILLER_12_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q net3278 VGND VPWR i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[138\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2582 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_99_126 VPWR VGND sg13g2_decap_8
XFILLER_5_583 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[110\]
+ net2997 i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y VPWR VGND i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_a21oi_1_A1_Y
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_o21ai_1_A1_Y
+ net3089 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_96_866 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[5\]_sg13g2_a22oi_1_A1 shift_reg_q\[5\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ net3053 net3044 net474 VPWR VGND sg13g2_a22oi_1
XFILLER_83_549 VPWR VGND sg13g2_decap_8
Xdata_pdata\[24\]_sg13g2_a21oi_1_A2 VGND VPWR data_pdata\[16\]_sg13g2_nor2b_1_B_N_Y
+ data_pdata\[24\]_sg13g2_a21oi_1_A2_Y data_pdata\[24\] net3159 sg13g2_a21oi_2
XFILLER_49_793 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nor2b_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y
+ net2925 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ net2923 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_76_590 VPWR VGND sg13g2_fill_2
XFILLER_48_281 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 net2761 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ net2519 VPWR VGND sg13g2_a22oi_1
XFILLER_64_774 VPWR VGND sg13g2_fill_1
XFILLER_36_465 VPWR VGND sg13g2_decap_4
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_36_498 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net3094 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[316\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_23_148 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2377
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[434\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2464 net2273 net2383 net1146 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net675 i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2372 net2738 i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y
+ net2569 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[482\]_sg13g2_nor3_1_A net1307 net2855 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[482\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_106_927 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1
+ net2579 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2
+ net2544 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A VGND VPWR
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 sg13g2_or2_1
XFILLER_59_524 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[435\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[435\]
+ net2999 i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_a21oi_1_A1_Y net2973 sg13g2_a21oi_1
XFILLER_87_888 VPWR VGND sg13g2_decap_8
XFILLER_101_698 VPWR VGND sg13g2_decap_4
XFILLER_98_1018 VPWR VGND sg13g2_decap_8
XFILLER_55_741 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[158\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_70_744 VPWR VGND sg13g2_fill_2
XFILLER_54_295 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2348
+ sg13g2_o21ai_1
XFILLER_35_1002 VPWR VGND sg13g2_fill_1
XFILLER_23_682 VPWR VGND sg13g2_fill_2
XFILLER_23_693 VPWR VGND sg13g2_decap_8
XFILLER_22_192 VPWR VGND sg13g2_decap_8
XFILLER_7_859 VPWR VGND sg13g2_fill_2
XFILLER_7_848 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[123\]
+ net2800 i_snitch.i_snitch_regfile.mem\[123\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xshift_reg_q\[5\]_sg13g2_nor2_1_A net474 net2730 shift_reg_q\[5\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xfanout3213 net3216 net3213 VPWR VGND sg13g2_buf_8
Xfanout3202 net3205 net3202 VPWR VGND sg13g2_buf_8
Xfanout3246 net3247 net3246 VPWR VGND sg13g2_buf_8
Xfanout3235 net3236 net3235 VPWR VGND sg13g2_buf_8
Xfanout2501 net2502 net2501 VPWR VGND sg13g2_buf_8
Xfanout3224 net3225 net3224 VPWR VGND sg13g2_buf_8
Xfanout2545 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y
+ net2545 VPWR VGND sg13g2_buf_8
XFILLER_78_800 VPWR VGND sg13g2_decap_4
Xfanout2523 net2529 net2523 VPWR VGND sg13g2_buf_8
Xfanout2534 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B_Y
+ net2534 VPWR VGND sg13g2_buf_8
Xfanout2512 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X
+ net2512 VPWR VGND sg13g2_buf_8
Xfanout3257 net3258 net3257 VPWR VGND sg13g2_buf_2
Xfanout3268 net3271 net3268 VPWR VGND sg13g2_buf_8
Xfanout3279 net3281 net3279 VPWR VGND sg13g2_buf_8
Xfanout2556 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y
+ net2556 VPWR VGND sg13g2_buf_8
Xfanout2578 net2579 net2578 VPWR VGND sg13g2_buf_8
Xfanout2567 net2568 net2567 VPWR VGND sg13g2_buf_8
Xuio_out_sg13g2_inv_1_Y_3 VPWR net9 uio_out_sg13g2_inv_1_Y_3_A VGND sg13g2_inv_1
Xfanout2589 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X
+ net2589 VPWR VGND sg13g2_buf_8
XFILLER_77_398 VPWR VGND sg13g2_fill_1
XFILLER_93_51 VPWR VGND sg13g2_fill_1
XFILLER_92_335 VPWR VGND sg13g2_fill_1
XFILLER_65_549 VPWR VGND sg13g2_fill_2
XFILLER_18_443 VPWR VGND sg13g2_decap_4
XFILLER_19_966 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_A1
+ net2308 i_snitch.pc_d\[21\] i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
XFILLER_73_571 VPWR VGND sg13g2_fill_2
XFILLER_73_560 VPWR VGND sg13g2_fill_1
XFILLER_45_240 VPWR VGND sg13g2_fill_1
XFILLER_18_476 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2374 net856 net2899 net2742 VPWR VGND sg13g2_a22oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C
+ net2641 i_snitch.i_snitch_regfile.mem\[470\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_60_265 VPWR VGND sg13g2_fill_2
XFILLER_60_254 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_40_clk clknet_5_11__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1
+ net2759 sg13g2_or2_1
Xstate_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net3053 cnt_q\[2\]_sg13g2_a22oi_1_B2_B1
+ state_sg13g2_dfrbpq_1_Q_D state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1 net2528 VPWR VGND sg13g2_xnor2_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2
+ net2512 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X VPWR
+ VGND sg13g2_and2_1
XFILLER_68_321 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[178\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_96_663 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2868
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_56_516 VPWR VGND sg13g2_fill_2
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
XFILLER_95_195 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2816 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_37_785 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B
+ net2517 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1 VPWR VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N
+ sg13g2_nand3b_1
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_24_435 VPWR VGND sg13g2_fill_2
XFILLER_36_284 VPWR VGND sg13g2_fill_2
XFILLER_11_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_31_clk clknet_5_14__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
Xdata_pdata\[0\]_sg13g2_mux2_1_A1 rsp_data_q\[0\] net684 net3051 data_pdata\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_32_490 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y net2956
+ i_snitch.i_snitch_regfile.mem\[282\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2961
+ i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[410\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
XFILLER_106_713 VPWR VGND sg13g2_decap_8
XFILLER_105_245 VPWR VGND sg13g2_decap_8
XFILLER_65_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_99_490 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_98_clk clknet_5_16__leaf_clk clknet_leaf_98_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[474\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[474\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net1099 net2460 net2255 VPWR VGND sg13g2_a22oi_1
XFILLER_75_803 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ net1227 VGND sg13g2_inv_1
XFILLER_102_996 VPWR VGND sg13g2_decap_8
XFILLER_47_538 VPWR VGND sg13g2_decap_4
XFILLER_74_346 VPWR VGND sg13g2_decap_4
XFILLER_28_752 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q
+ net3195 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[16\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
XFILLER_15_402 VPWR VGND sg13g2_fill_1
XFILLER_43_722 VPWR VGND sg13g2_decap_8
XFILLER_16_936 VPWR VGND sg13g2_decap_8
XFILLER_43_766 VPWR VGND sg13g2_decap_4
XFILLER_15_468 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_o21ai_1_A1_B1
+ i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_o21ai_1_A1_Y VGND sg13g2_inv_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_Y
+ i_req_arb.data_i\[37\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C
+ net2533 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A
+ VPWR VGND sg13g2_nor4_1
Xclkbuf_leaf_22_clk clknet_5_14__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_8_49 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ net2573 net2538 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_a21o_1
XFILLER_6_133 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_o21ai_1_A1 net2970 VPWR i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[365\] net2804 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q net3293 VGND VPWR i_snitch.i_snitch_regfile.mem\[198\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[198\] clknet_leaf_78_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[504\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[504\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_98_906 VPWR VGND sg13g2_decap_8
Xfanout3021 net3023 net3021 VPWR VGND sg13g2_buf_8
Xfanout3010 net3011 net3010 VPWR VGND sg13g2_buf_8
Xfanout3032 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net3032 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y
+ net439 VGND sg13g2_inv_1
Xfanout3043 net3044 net3043 VPWR VGND sg13g2_buf_8
Xcnt_q\[2\]_sg13g2_a21oi_1_B1 VGND VPWR cnt_q\[1\] cnt_q\[0\] cnt_q\[2\]_sg13g2_a21oi_1_B1_Y
+ net448 sg13g2_a21oi_1
Xfanout3054 net3055 net3054 VPWR VGND sg13g2_buf_1
Xfanout2320 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2320 VPWR VGND sg13g2_buf_8
Xfanout3076 net3077 net3076 VPWR VGND sg13g2_buf_8
Xfanout3065 net3067 net3065 VPWR VGND sg13g2_buf_8
Xfanout3087 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ net3087 VPWR VGND sg13g2_buf_8
Xfanout3098 net3099 net3098 VPWR VGND sg13g2_buf_8
Xfanout2353 net2354 net2353 VPWR VGND sg13g2_buf_8
Xfanout2342 net2346 net2342 VPWR VGND sg13g2_buf_8
Xfanout2331 net2333 net2331 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ sg13g2_nand2b_2
Xfanout2375 net2376 net2375 VPWR VGND sg13g2_buf_8
Xfanout2386 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2386 VPWR VGND sg13g2_buf_8
Xfanout2364 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ net2364 VPWR VGND sg13g2_buf_2
Xclkbuf_leaf_89_clk clknet_5_21__leaf_clk clknet_leaf_89_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[46\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_78_696 VPWR VGND sg13g2_decap_8
XFILLER_66_836 VPWR VGND sg13g2_decap_4
XFILLER_38_527 VPWR VGND sg13g2_decap_8
Xfanout2397 net2398 net2397 VPWR VGND sg13g2_buf_8
XFILLER_92_132 VPWR VGND sg13g2_fill_2
XFILLER_66_869 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2482 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2532 VPWR VGND sg13g2_a22oi_1
XFILLER_65_335 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21o_1_X
+ net2491 net666 net2429 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_a21o_1
XFILLER_80_327 VPWR VGND sg13g2_fill_1
XFILLER_46_571 VPWR VGND sg13g2_decap_8
XFILLER_61_552 VPWR VGND sg13g2_fill_2
XFILLER_22_917 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y net2841 i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_34_799 VPWR VGND sg13g2_fill_2
XFILLER_105_1022 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_5_6__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2874
+ i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xdata_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A_Y net2842 i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_30_972 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[494\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2368 net952 net2688 net2857 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2661 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A net1358 net2868 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C
+ i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[258\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[258\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[258\] VGND sg13g2_inv_1
XFILLER_88_416 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q
+ net3203 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_102_259 VPWR VGND sg13g2_decap_8
XFILLER_97_950 VPWR VGND sg13g2_decap_8
XFILLER_69_652 VPWR VGND sg13g2_decap_8
XFILLER_68_140 VPWR VGND sg13g2_decap_4
XFILLER_57_825 VPWR VGND sg13g2_fill_1
XFILLER_68_195 VPWR VGND sg13g2_fill_1
XFILLER_57_869 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2771
+ net2673 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_Y
+ VPWR VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[354\]_sg13g2_nor3_1_A net1334 net2879 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_52_552 VPWR VGND sg13g2_fill_2
XFILLER_24_232 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_A1
+ net2304 i_snitch.pc_d\[28\] i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2430 net2267 net2316 net1268 VPWR VGND sg13g2_a22oi_1
XFILLER_21_983 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[66\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[66\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[66\] clknet_leaf_108_clk sg13g2_dfrbpq_1
XFILLER_106_565 VPWR VGND sg13g2_decap_8
XFILLER_79_416 VPWR VGND sg13g2_decap_8
XFILLER_0_821 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[314\]
+ net3000 i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_a21oi_1_A1_Y net2976 sg13g2_a21oi_1
XFILLER_88_994 VPWR VGND sg13g2_decap_8
XFILLER_59_140 VPWR VGND sg13g2_fill_1
XFILLER_58_87 VPWR VGND sg13g2_fill_1
XFILLER_48_814 VPWR VGND sg13g2_decap_8
XFILLER_0_898 VPWR VGND sg13g2_decap_8
XFILLER_102_793 VPWR VGND sg13g2_decap_8
XFILLER_75_688 VPWR VGND sg13g2_decap_4
Xi_snitch.inst_addr_o\[18\]_sg13g2_inv_1_A i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1
+ net1355 VPWR VGND sg13g2_inv_2
Xdata_pdata\[8\]_sg13g2_nand2b_1_B data_pdata\[8\]_sg13g2_nand2b_1_B_Y data_pdata\[8\]
+ net3159 VPWR VGND sg13g2_nand2b_1
XFILLER_47_357 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2294 net1347 net2491 net1212 VPWR VGND sg13g2_a22oi_1
XFILLER_16_744 VPWR VGND sg13g2_decap_8
Xdata_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[8\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[24\]_sg13g2_nand2b_1_B_Y net3152 data_pdata\[16\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[8\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
XFILLER_43_596 VPWR VGND sg13g2_decap_8
XFILLER_30_213 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ VGND net2712 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[388\] VGND sg13g2_inv_1
Xhold409 i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A
+ VPWR VGND net441 sg13g2_dlygate4sd3_1
Xdata_pdata\[7\]_sg13g2_mux2_1_A1 rsp_data_q\[7\] net681 net3051 data_pdata\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_976 VPWR VGND sg13g2_decap_8
Xdata_pdata\[7\]_sg13g2_dfrbpq_1_Q net3228 VGND VPWR net682 data_pdata\[7\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_3_681 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2898 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2456 VPWR VGND sg13g2_nand2_1
XFILLER_86_909 VPWR VGND sg13g2_decap_8
XFILLER_31_4 VPWR VGND sg13g2_fill_1
XFILLER_94_931 VPWR VGND sg13g2_decap_8
XFILLER_79_972 VPWR VGND sg13g2_decap_8
Xhold1109 i_snitch.i_snitch_regfile.mem\[373\] VPWR VGND net1141 sg13g2_dlygate4sd3_1
Xcnt_q\[2\]_sg13g2_a22oi_1_B2_B1_sg13g2_nand2_1_Y cnt_q\[2\]_sg13g2_a22oi_1_B2_B1
+ net1 strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B1 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_2_clk clknet_5_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_65_110 VPWR VGND sg13g2_decap_4
XFILLER_93_463 VPWR VGND sg13g2_fill_1
XFILLER_93_452 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2405 net976 net2689 net2798 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y_sg13g2_nor2b_1_A
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2b_2
XFILLER_65_176 VPWR VGND sg13g2_fill_2
XFILLER_53_338 VPWR VGND sg13g2_fill_2
XFILLER_0_1003 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q net3320 VGND VPWR i_snitch.i_snitch_regfile.mem\[86\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[86\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_80_168 VPWR VGND sg13g2_fill_1
XFILLER_55_1027 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]
+ net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2 i_snitch.inst_addr_o\[11\] i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2542 VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ VGND net2750 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ sg13g2_o21ai_1
Xhold921 i_snitch.i_snitch_regfile.mem\[168\] VPWR VGND net953 sg13g2_dlygate4sd3_1
Xhold910 data_pdata\[27\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net942 sg13g2_dlygate4sd3_1
Xhold943 i_snitch.i_snitch_regfile.mem\[401\] VPWR VGND net975 sg13g2_dlygate4sd3_1
Xhold954 i_snitch.i_snitch_regfile.mem\[370\] VPWR VGND net986 sg13g2_dlygate4sd3_1
Xhold932 i_snitch.i_snitch_regfile.mem\[350\] VPWR VGND net964 sg13g2_dlygate4sd3_1
Xhold987 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net1019 sg13g2_dlygate4sd3_1
Xhold998 i_snitch.i_snitch_regfile.mem\[271\] VPWR VGND net1030 sg13g2_dlygate4sd3_1
XFILLER_1_629 VPWR VGND sg13g2_decap_8
Xhold976 i_snitch.i_snitch_regfile.mem\[455\] VPWR VGND net1008 sg13g2_dlygate4sd3_1
Xhold965 i_snitch.i_snitch_regfile.mem\[330\] VPWR VGND net997 sg13g2_dlygate4sd3_1
XFILLER_103_557 VPWR VGND sg13g2_decap_8
XFILLER_89_758 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[190\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2774
+ net2649 VPWR VGND sg13g2_nand2_1
Xi_snitch.gpr_waddr\[7\]_sg13g2_nor2_1_A i_snitch.gpr_waddr\[7\] i_snitch.gpr_waddr\[6\]
+ i_snitch.gpr_waddr\[7\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_85_920 VPWR VGND sg13g2_decap_8
XFILLER_57_600 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_mux2_1_A1
+ net537 net619 net2617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_28_46 VPWR VGND sg13g2_fill_2
XFILLER_29_324 VPWR VGND sg13g2_fill_2
XFILLER_85_997 VPWR VGND sg13g2_decap_8
XFILLER_84_474 VPWR VGND sg13g2_fill_2
XFILLER_84_463 VPWR VGND sg13g2_decap_8
XFILLER_84_452 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_44_338 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ VGND net2712 i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
XFILLER_25_530 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y
+ net55 VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B
+ VGND net2566 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ sg13g2_a21oi_2
XFILLER_44_56 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR net58 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_inv_1_A_Y
+ net2622 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_12_213 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2431
+ net2287 VPWR VGND sg13g2_nand2_1
XFILLER_40_566 VPWR VGND sg13g2_decap_8
XFILLER_100_84 VPWR VGND sg13g2_decap_8
Xi_req_register.data_o\[39\]_sg13g2_o21ai_1_Y i_req_register.data_o\[39\]_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.data_o\[39\] VGND net3173 i_req_register.data_o\[39\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2837 i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_40_599 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y net2918 i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net3092 sg13g2_a21oi_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1
+ VPWR VGND sg13g2_nor2_1
XFILLER_5_935 VPWR VGND sg13g2_decap_8
Xdata_pdata\[19\]_sg13g2_mux2_1_A0 data_pdata\[19\] data_pdata\[27\] net3158 data_pdata\[19\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_5_39 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.pc_d\[1\]
+ VGND net2301 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[398\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2468 VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2
+ net2506 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_95_717 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ net2547 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_xor2_1
XFILLER_0_695 VPWR VGND sg13g2_decap_8
XFILLER_91_912 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ net69 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_76_997 VPWR VGND sg13g2_decap_8
XFILLER_90_422 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A
+ VGND VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A sg13g2_or2_1
XFILLER_62_113 VPWR VGND sg13g2_fill_2
XFILLER_91_989 VPWR VGND sg13g2_decap_8
XFILLER_90_466 VPWR VGND sg13g2_decap_8
XFILLER_90_433 VPWR VGND sg13g2_decap_8
XFILLER_16_541 VPWR VGND sg13g2_decap_8
XFILLER_18_90 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] net571 net2616
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ net1139 net1093 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_102_1003 VPWR VGND sg13g2_decap_8
XFILLER_7_294 VPWR VGND sg13g2_fill_2
XFILLER_98_533 VPWR VGND sg13g2_fill_1
XFILLER_4_990 VPWR VGND sg13g2_decap_8
XFILLER_59_909 VPWR VGND sg13g2_decap_8
XFILLER_100_527 VPWR VGND sg13g2_decap_8
XFILLER_100_516 VPWR VGND sg13g2_fill_1
XFILLER_61_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C net414
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C net2762 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ net45 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_67_964 VPWR VGND sg13g2_decap_8
XFILLER_94_794 VPWR VGND sg13g2_decap_4
XFILLER_82_923 VPWR VGND sg13g2_decap_8
Xi_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y VGND VPWR i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1
+ net70 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ sg13g2_nand2b_2
XFILLER_66_496 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_dfrbpq_1_Q
+ net3192 VGND VPWR net663 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
XFILLER_93_293 VPWR VGND sg13g2_decap_4
XFILLER_53_146 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_and2_1
XFILLER_50_864 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net1141 net2469 net2269 VPWR VGND sg13g2_a22oi_1
XFILLER_5_209 VPWR VGND sg13g2_decap_4
XFILLER_100_7 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2580 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xhold740 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] VPWR
+ VGND net772 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold751 i_snitch.i_snitch_regfile.mem\[224\] VPWR VGND net783 sg13g2_dlygate4sd3_1
Xhold762 i_snitch.i_snitch_regfile.mem\[73\] VPWR VGND net794 sg13g2_dlygate4sd3_1
XFILLER_1_415 VPWR VGND sg13g2_decap_4
Xfanout2919 net81 net2919 VPWR VGND sg13g2_buf_8
Xhold773 i_snitch.i_snitch_regfile.mem\[429\] VPWR VGND net805 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[226\]_sg13g2_nor3_1_A net1357 net2872 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[226\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xfanout2908 data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y net2908 VPWR VGND
+ sg13g2_buf_8
XFILLER_104_844 VPWR VGND sg13g2_decap_8
XFILLER_103_343 VPWR VGND sg13g2_decap_8
Xhold795 i_snitch.i_snitch_regfile.mem\[408\] VPWR VGND net827 sg13g2_dlygate4sd3_1
Xhold784 i_snitch.i_snitch_regfile.mem\[424\] VPWR VGND net816 sg13g2_dlygate4sd3_1
XFILLER_77_728 VPWR VGND sg13g2_fill_2
XFILLER_49_408 VPWR VGND sg13g2_decap_8
XFILLER_55_11 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[508\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2458 net2247 net2369 net1324 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_45_647 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A VPWR
+ VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q net3208 VGND VPWR i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[403\] clknet_leaf_120_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]
+ net3164 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_41_875 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[509\]
+ net3127 i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1
+ net2923 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2
+ sg13g2_a221oi_1
XFILLER_5_721 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2377
+ sg13g2_o21ai_1
XFILLER_4_297 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_dfrbpq_1_Q
+ net3195 VGND VPWR net425 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
Xi_snitch.sb_q\[9\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.sb_d\[9\] i_snitch.sb_q\[9\]
+ clknet_leaf_106_clk sg13g2_dfrbpq_1
XFILLER_96_84 VPWR VGND sg13g2_decap_8
XFILLER_95_558 VPWR VGND sg13g2_decap_4
XFILLER_95_525 VPWR VGND sg13g2_fill_1
XFILLER_1_993 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D_sg13g2_and2_1_X
+ net3147 net3073 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D
+ VPWR VGND sg13g2_and2_1
XFILLER_91_731 VPWR VGND sg13g2_fill_2
XFILLER_64_945 VPWR VGND sg13g2_decap_8
XFILLER_64_956 VPWR VGND sg13g2_fill_1
XFILLER_63_455 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[393\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[393\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2388 net800 net2685 net3039 VPWR VGND sg13g2_a22oi_1
XFILLER_17_850 VPWR VGND sg13g2_fill_1
XFILLER_91_797 VPWR VGND sg13g2_decap_8
XFILLER_91_1024 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[112\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2759 net2307
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2520 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[394\]
+ net3027 i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[426\]_sg13g2_a21o_1_A1_X
+ sg13g2_a21oi_1
XFILLER_99_853 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[7\] net772 net2914 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[284\] net2814 sg13g2_o21ai_1
XFILLER_101_847 VPWR VGND sg13g2_decap_8
XFILLER_100_324 VPWR VGND sg13g2_decap_8
XFILLER_86_525 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[423\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[423\] clknet_leaf_118_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]
+ net3167 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_86_569 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2363
+ sg13g2_o21ai_1
XFILLER_94_580 VPWR VGND sg13g2_decap_4
Xrebuffer21 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ net53 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[212\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[212\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net718 net2671 net2791 VPWR VGND sg13g2_a22oi_1
Xrebuffer10 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ net42 VPWR VGND sg13g2_buf_1
XFILLER_94_591 VPWR VGND sg13g2_decap_4
Xrebuffer43 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y
+ net75 VPWR VGND sg13g2_buf_1
Xrebuffer54 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y
+ net86 VPWR VGND sg13g2_buf_1
XFILLER_81_230 VPWR VGND sg13g2_decap_4
Xrebuffer32 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y
+ net64 VPWR VGND sg13g2_buf_1
Xrebuffer87 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D
+ net119 VPWR VGND sg13g2_buf_1
Xrebuffer76 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y
+ net108 VPWR VGND sg13g2_buf_1
Xrebuffer65 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X
+ net97 VPWR VGND sg13g2_buf_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y
+ net3175 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_25_69 VPWR VGND sg13g2_fill_2
XFILLER_35_680 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\] net594 net2623
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[29\]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A i_snitch.pc_d\[26\]_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[16\]_sg13g2_a221oi_1_A2_Y i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D_Y
+ i_snitch.pc_d\[29\]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A_Y VPWR VGND i_snitch.pc_d\[29\]_sg13g2_nand2_1_B_Y
+ sg13g2_nand4_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2771
+ i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y
+ net2613 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ VPWR VGND sg13g2_nor4_1
XFILLER_41_68 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y
+ VGND VPWR net89 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y
+ sg13g2_nand2b_2
Xfanout2705 net2708 net2705 VPWR VGND sg13g2_buf_8
Xfanout2716 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y
+ net2716 VPWR VGND sg13g2_buf_8
Xfanout2727 net2729 net2727 VPWR VGND sg13g2_buf_8
Xhold570 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net602 sg13g2_dlygate4sd3_1
Xhold581 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net613 sg13g2_dlygate4sd3_1
XFILLER_103_140 VPWR VGND sg13g2_decap_8
Xfanout2749 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1_X
+ net2749 VPWR VGND sg13g2_buf_8
Xhold592 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net624 sg13g2_dlygate4sd3_1
Xfanout2738 net2740 net2738 VPWR VGND sg13g2_buf_8
XFILLER_2_768 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[103\]
+ net2947 sg13g2_o21ai_1
XFILLER_2_18 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2485 i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2471 net2879 i_snitch.i_snitch_regfile.mem\[354\]_sg13g2_dfrbpq_1_Q_D net2912
+ sg13g2_a221oi_1
XFILLER_77_558 VPWR VGND sg13g2_fill_1
XFILLER_85_580 VPWR VGND sg13g2_fill_2
XFILLER_17_102 VPWR VGND sg13g2_fill_2
XFILLER_18_603 VPWR VGND sg13g2_fill_2
Xhold1270 i_snitch.i_snitch_regfile.mem\[106\] VPWR VGND net1302 sg13g2_dlygate4sd3_1
XFILLER_57_282 VPWR VGND sg13g2_decap_8
XFILLER_45_433 VPWR VGND sg13g2_fill_2
Xhold1292 i_snitch.i_snitch_regfile.mem\[508\] VPWR VGND net1324 sg13g2_dlygate4sd3_1
Xhold1281 i_snitch.i_snitch_regfile.mem\[484\] VPWR VGND net1313 sg13g2_dlygate4sd3_1
XFILLER_26_691 VPWR VGND sg13g2_decap_4
Xheichips25_snitch_wrapper_25 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_25_190 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1
+ VPWR VGND net2933 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ net3088 sg13g2_a221oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y
+ sg13g2_a21oi_2
XFILLER_41_683 VPWR VGND sg13g2_fill_2
XFILLER_9_345 VPWR VGND sg13g2_fill_2
XFILLER_9_378 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nand2b_1_A_N
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y_B1
+ net2707 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[443\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[443\] clknet_leaf_119_clk sg13g2_dfrbpq_1
XFILLER_99_105 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1
+ net531 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[232\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[232\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2331 net1137 net2643 net2875 VPWR VGND sg13g2_a22oi_1
XFILLER_96_845 VPWR VGND sg13g2_decap_8
XFILLER_95_300 VPWR VGND sg13g2_fill_2
XFILLER_1_790 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[3\]_sg13g2_nor2_1_A net459 net2727 strb_reg_q\[3\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_91_550 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[439\]_sg13g2_o21ai_1_A1 net3096 VPWR i_snitch.i_snitch_regfile.mem\[439\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[439\] net2812 sg13g2_o21ai_1
XFILLER_51_403 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[19\]_sg13g2_nor2_1_A net498 net2733 shift_reg_q\[19\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_36_488 VPWR VGND sg13g2_decap_4
XFILLER_17_680 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q
+ net3235 VGND VPWR net1043 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
XFILLER_51_469 VPWR VGND sg13g2_fill_2
XFILLER_16_190 VPWR VGND sg13g2_decap_4
XFILLER_32_661 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2614 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_20_878 VPWR VGND sg13g2_decap_8
XFILLER_106_906 VPWR VGND sg13g2_decap_8
XFILLER_105_427 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_nand2b_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2762 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
Xrsp_data_q\[24\]_sg13g2_dfrbpq_1_Q net3238 VGND VPWR rsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[24\] clknet_leaf_34_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[440\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2380
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2420 sg13g2_a21oi_1
XFILLER_101_633 VPWR VGND sg13g2_fill_2
XFILLER_98_182 VPWR VGND sg13g2_fill_1
XFILLER_87_867 VPWR VGND sg13g2_decap_8
XFILLER_59_569 VPWR VGND sg13g2_decap_8
XFILLER_100_154 VPWR VGND sg13g2_decap_8
XFILLER_46_208 VPWR VGND sg13g2_decap_8
XFILLER_100_198 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y
+ net2848 net52 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_nor2_2
XFILLER_55_731 VPWR VGND sg13g2_fill_1
XFILLER_55_797 VPWR VGND sg13g2_fill_1
XFILLER_54_274 VPWR VGND sg13g2_decap_8
XFILLER_15_639 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[183\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2341
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[463\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[463\] clknet_leaf_81_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[252\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[252\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net1024 net2437 net2246 VPWR VGND sg13g2_a22oi_1
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1 net545 i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xfanout3203 net3205 net3203 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[430\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net455 net2381 VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2479 net2416 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2499 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y
+ sg13g2_a221oi_1
Xfanout3247 net3248 net3247 VPWR VGND sg13g2_buf_8
Xfanout3236 net3249 net3236 VPWR VGND sg13g2_buf_8
Xfanout2502 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A_Y
+ net2502 VPWR VGND sg13g2_buf_8
Xfanout3214 net3216 net3214 VPWR VGND sg13g2_buf_8
Xfanout3225 net3226 net3225 VPWR VGND sg13g2_buf_8
XFILLER_81_1012 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y VPWR i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_A1
+ net1242 VGND sg13g2_inv_1
Xfanout2524 net2529 net2524 VPWR VGND sg13g2_buf_2
Xfanout2535 net2535 net2536 VPWR VGND sg13g2_buf_16
Xfanout3258 net3259 net3258 VPWR VGND sg13g2_buf_8
Xfanout3269 net3271 net3269 VPWR VGND sg13g2_buf_8
Xfanout2513 net2514 net2513 VPWR VGND sg13g2_buf_8
XFILLER_105_994 VPWR VGND sg13g2_decap_8
Xfanout2557 net2559 net2557 VPWR VGND sg13g2_buf_8
Xfanout2546 net2547 net2546 VPWR VGND sg13g2_buf_8
XFILLER_89_160 VPWR VGND sg13g2_fill_1
Xfanout2568 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1_Y
+ net2568 VPWR VGND sg13g2_buf_8
XFILLER_78_856 VPWR VGND sg13g2_decap_8
Xfanout2579 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y
+ net2579 VPWR VGND sg13g2_buf_8
XFILLER_78_867 VPWR VGND sg13g2_fill_2
XFILLER_65_506 VPWR VGND sg13g2_fill_2
XFILLER_65_528 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR net652 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_37_208 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1
+ net2705 i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_46_753 VPWR VGND sg13g2_fill_1
XFILLER_19_945 VPWR VGND sg13g2_fill_2
XFILLER_46_786 VPWR VGND sg13g2_fill_2
XFILLER_19_978 VPWR VGND sg13g2_fill_2
XFILLER_34_904 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2601 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_61_723 VPWR VGND sg13g2_fill_1
XFILLER_60_222 VPWR VGND sg13g2_fill_1
XFILLER_45_285 VPWR VGND sg13g2_decap_4
XFILLER_33_425 VPWR VGND sg13g2_fill_2
XFILLER_61_767 VPWR VGND sg13g2_fill_2
XFILLER_33_458 VPWR VGND sg13g2_fill_1
Xrebuffer1 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D_Y
+ net33 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A_Y net2985 i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net3028 sg13g2_a21oi_1
XFILLER_68_300 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0 net3129 i_snitch.i_snitch_regfile.mem\[146\]
+ i_snitch.i_snitch_regfile.mem\[178\] i_snitch.i_snitch_regfile.mem\[210\] i_snitch.i_snitch_regfile.mem\[242\]
+ net3108 i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[483\] clknet_leaf_100_clk sg13g2_dfrbpq_1
XFILLER_28_208 VPWR VGND sg13g2_decap_8
XFILLER_28_219 VPWR VGND sg13g2_fill_2
Xdata_pdata\[26\]_sg13g2_nand2b_1_B data_pdata\[26\]_sg13g2_nand2b_1_B_Y data_pdata\[26\]
+ net3156 VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net1229 net2434 net2263 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2530 i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_64_550 VPWR VGND sg13g2_decap_4
XFILLER_92_892 VPWR VGND sg13g2_decap_8
XFILLER_51_200 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2935 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_25_959 VPWR VGND sg13g2_decap_8
XFILLER_51_255 VPWR VGND sg13g2_decap_4
XFILLER_51_233 VPWR VGND sg13g2_fill_2
Xcnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D VGND cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A
+ cnt_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_51_277 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1 net2967 VPWR i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[479\] i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_A2
+ sg13g2_o21ai_1
XFILLER_22_37 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.sb_q\[9\] net3008 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1
+ net2980 sg13g2_a21oi_1
XFILLER_105_224 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[407\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net898 net2647 net3041 VPWR VGND sg13g2_a22oi_1
XFILLER_3_329 VPWR VGND sg13g2_fill_1
Xdata_pdata\[25\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net946 data_pdata\[25\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
XFILLER_87_642 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q net3292 VGND VPWR i_snitch.i_snitch_regfile.mem\[302\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[302\] clknet_leaf_85_clk sg13g2_dfrbpq_1
XFILLER_102_975 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_A1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A
+ VGND sg13g2_inv_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2_sg13g2_nor2b_1_Y
+ net3144 net3142 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2
+ VPWR VGND sg13g2_nor2b_2
XFILLER_75_815 VPWR VGND sg13g2_decap_8
XFILLER_16_904 VPWR VGND sg13g2_decap_8
XFILLER_103_84 VPWR VGND sg13g2_decap_8
XFILLER_82_380 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[408\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[408\]
+ net3030 i_snitch.i_snitch_regfile.mem\[408\]_sg13g2_a21oi_1_A1_Y net2993 sg13g2_a21oi_1
XFILLER_55_583 VPWR VGND sg13g2_decap_4
XFILLER_27_263 VPWR VGND sg13g2_decap_8
XFILLER_70_542 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[105\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[105\] VGND sg13g2_inv_1
XFILLER_30_417 VPWR VGND sg13g2_fill_1
XFILLER_31_929 VPWR VGND sg13g2_decap_4
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_fill_1
XFILLER_10_152 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_mux2_1_A1 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[23\]
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_A1 i_snitch.pc_d\[23\]_sg13g2_mux2_1_A1_X VPWR
+ VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A_sg13g2_nor2_1_Y
+ net49 net2500 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ VPWR VGND sg13g2_nor2_2
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_6_167 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ net2613 VPWR VGND sg13g2_a22oi_1
XFILLER_88_30 VPWR VGND sg13g2_decap_4
Xfanout3022 net3023 net3022 VPWR VGND sg13g2_buf_8
Xfanout3000 net3003 net3000 VPWR VGND sg13g2_buf_8
Xfanout3011 net3025 net3011 VPWR VGND sg13g2_buf_8
Xfanout3033 net3034 net3033 VPWR VGND sg13g2_buf_8
Xfanout2310 net106 net2310 VPWR VGND sg13g2_buf_2
Xfanout3055 state_sg13g2_inv_1_A_Y net3055 VPWR VGND sg13g2_buf_8
Xfanout3044 net3045 net3044 VPWR VGND sg13g2_buf_8
XFILLER_105_791 VPWR VGND sg13g2_decap_8
XFILLER_97_439 VPWR VGND sg13g2_fill_1
Xfanout3077 net3078 net3077 VPWR VGND sg13g2_buf_8
Xfanout3066 net3067 net3066 VPWR VGND sg13g2_buf_8
XFILLER_69_119 VPWR VGND sg13g2_fill_1
Xfanout3088 net3090 net3088 VPWR VGND sg13g2_buf_8
Xfanout2321 net2322 net2321 VPWR VGND sg13g2_buf_8
Xfanout2343 net2346 net2343 VPWR VGND sg13g2_buf_8
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_2_384 VPWR VGND sg13g2_fill_1
Xfanout2332 net2333 net2332 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[31\] net831 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0 net3122 i_snitch.i_snitch_regfile.mem\[384\]
+ i_snitch.i_snitch_regfile.mem\[416\] i_snitch.i_snitch_regfile.mem\[448\] i_snitch.i_snitch_regfile.mem\[480\]
+ net3104 i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xfanout2365 net2366 net2365 VPWR VGND sg13g2_buf_8
Xfanout3099 net3102 net3099 VPWR VGND sg13g2_buf_8
Xfanout2354 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2354 VPWR VGND sg13g2_buf_8
Xfanout2387 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2387 VPWR VGND sg13g2_buf_8
Xfanout2376 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2376 VPWR VGND sg13g2_buf_8
Xdata_pdata\[17\]_sg13g2_a21oi_1_A2 VGND VPWR net3155 data_pdata\[17\] data_pdata\[17\]_sg13g2_a21oi_1_A2_Y
+ net3149 sg13g2_a21oi_1
Xfanout2398 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2398 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR
+ net2486 net2501 i_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D i_snitch.i_snitch_lsu.metadata_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_92_144 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[499\]_sg13g2_o21ai_1_A1 net2961 VPWR i_snitch.i_snitch_regfile.mem\[499\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[499\] net2800 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[293\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[293\]
+ net3001 i_snitch.i_snitch_regfile.mem\[293\]_sg13g2_a21oi_1_A1_Y net2975 sg13g2_a21oi_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2603 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_18_1020 VPWR VGND sg13g2_decap_8
XFILLER_105_1001 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ net2927 net2744 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net1068 net2679 net2863 VPWR VGND sg13g2_a22oi_1
Xdata_pdata\[12\]_sg13g2_mux2_1_A1 rsp_data_q\[12\] net901 net3051 data_pdata\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR
+ VGND net2833 net2639 i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y net2954
+ i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[322\] clknet_leaf_109_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2412 net843 net2678 net2871 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3168 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A_Y
+ strb_reg_q\[2\]_sg13g2_a21oi_1_A1_B1 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
Xshift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[35\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y
+ VPWR shift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 VGND net3165 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]
+ sg13g2_o21ai_1
XFILLER_102_238 VPWR VGND sg13g2_decap_8
XFILLER_71_306 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[10\]_sg13g2_a22oi_1_A1 shift_reg_q\[10\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 net468 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[318\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[318\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[318\] net2812 sg13g2_o21ai_1
XFILLER_83_199 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2416 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_52_542 VPWR VGND sg13g2_fill_1
XFILLER_13_929 VPWR VGND sg13g2_fill_2
XFILLER_25_778 VPWR VGND sg13g2_decap_8
XFILLER_12_439 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_B1
+ net1074 net2304 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2590 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[479\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_106_544 VPWR VGND sg13g2_decap_4
XFILLER_58_11 VPWR VGND sg13g2_decap_8
XFILLER_0_800 VPWR VGND sg13g2_decap_8
Xdata_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2 data_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ net3070 net2714 data_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_88_973 VPWR VGND sg13g2_decap_8
XFILLER_58_99 VPWR VGND sg13g2_fill_1
XFILLER_0_877 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[447\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2382 net933 net2646 net2863 VPWR VGND sg13g2_a22oi_1
XFILLER_62_306 VPWR VGND sg13g2_decap_4
XFILLER_62_339 VPWR VGND sg13g2_fill_2
XFILLER_15_211 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[342\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_43_542 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[115\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2866
+ net2674 VPWR VGND sg13g2_nand2_1
XFILLER_16_767 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q
+ net3242 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_43_586 VPWR VGND sg13g2_decap_4
XFILLER_43_575 VPWR VGND sg13g2_fill_1
XFILLER_15_255 VPWR VGND sg13g2_decap_4
XFILLER_30_203 VPWR VGND sg13g2_fill_1
XFILLER_12_984 VPWR VGND sg13g2_decap_4
Xi_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q net3251 VGND VPWR i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.gpr_waddr\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[219\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2788
+ net2657 VPWR VGND sg13g2_nand2_1
XFILLER_99_84 VPWR VGND sg13g2_decap_8
XFILLER_98_715 VPWR VGND sg13g2_decap_8
XFILLER_98_726 VPWR VGND sg13g2_fill_1
XFILLER_3_660 VPWR VGND sg13g2_decap_8
XFILLER_79_951 VPWR VGND sg13g2_decap_8
XFILLER_94_910 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y net3017 sg13g2_o21ai_1
XFILLER_78_494 VPWR VGND sg13g2_fill_1
XFILLER_94_987 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2567 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_2
XFILLER_66_689 VPWR VGND sg13g2_fill_1
XFILLER_65_144 VPWR VGND sg13g2_fill_2
XFILLER_65_133 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[99\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_nor3_1_A_Y net2448 net2866 i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_dfrbpq_1_Q_D
+ net2909 sg13g2_a221oi_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2695 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ net2540 sg13g2_a21oi_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_xor2_1
XFILLER_94_1022 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2552 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y
+ sg13g2_a21oi_1
XFILLER_62_862 VPWR VGND sg13g2_fill_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_22_726 VPWR VGND sg13g2_fill_2
XFILLER_34_575 VPWR VGND sg13g2_fill_2
XFILLER_22_748 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_B i_snitch.inst_addr_o\[21\]
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_B1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1
+ net2748 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
Xhold922 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\] VPWR
+ VGND net954 sg13g2_dlygate4sd3_1
Xhold900 i_snitch.i_snitch_regfile.mem\[477\] VPWR VGND net932 sg13g2_dlygate4sd3_1
Xhold911 i_snitch.i_snitch_regfile.mem\[469\] VPWR VGND net943 sg13g2_dlygate4sd3_1
XFILLER_89_715 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net1159 net2460 net2270 VPWR VGND sg13g2_a22oi_1
XFILLER_1_608 VPWR VGND sg13g2_decap_8
Xhold955 i_snitch.i_snitch_regfile.mem\[71\] VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold944 i_snitch.i_snitch_regfile.mem\[333\] VPWR VGND net976 sg13g2_dlygate4sd3_1
Xhold933 i_snitch.i_snitch_regfile.mem\[134\] VPWR VGND net965 sg13g2_dlygate4sd3_1
XFILLER_103_525 VPWR VGND sg13g2_fill_1
Xhold966 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\] VPWR
+ VGND net998 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2889
+ net2675 VPWR VGND sg13g2_nand2_1
Xhold977 i_snitch.i_snitch_regfile.mem\[154\] VPWR VGND net1009 sg13g2_dlygate4sd3_1
Xhold988 i_snitch.i_snitch_regfile.mem\[266\] VPWR VGND net1020 sg13g2_dlygate4sd3_1
Xshift_reg_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2734 shift_reg_q\[27\]_sg13g2_a22oi_1_A1_Y
+ shift_reg_q\[23\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[23\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
Xhold999 i_snitch.i_snitch_regfile.mem\[359\] VPWR VGND net1031 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_or2_1_X VGND VPWR
+ i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q net3270 VGND VPWR i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[362\] clknet_leaf_102_clk sg13g2_dfrbpq_1
XFILLER_96_291 VPWR VGND sg13g2_fill_1
XFILLER_56_111 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1 VPWR VGND net3100 net2821
+ i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_mux2_1_A0_X i_snitch.i_snitch_regfile.mem\[57\]
+ i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1_Y net2824 sg13g2_a221oi_1
XFILLER_85_976 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2350 net851 net2648 net2888 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1322 net2495 net1177 VPWR VGND sg13g2_a22oi_1
XFILLER_40_501 VPWR VGND sg13g2_decap_8
XFILLER_40_545 VPWR VGND sg13g2_fill_1
XFILLER_100_63 VPWR VGND sg13g2_decap_8
Xdata_pdata\[2\]_sg13g2_nor2_1_B net3157 data_pdata\[2\] data_pdata\[2\]_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_5_914 VPWR VGND sg13g2_decap_8
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
Xdata_pdata\[19\]_sg13g2_mux2_1_A1 rsp_data_q\[19\] net754 net3049 data_pdata\[19\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_69_21 VPWR VGND sg13g2_fill_1
XFILLER_106_385 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[22\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[22\]
+ i_snitch.inst_addr_o\[22\] clknet_leaf_57_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q net3215 VGND VPWR i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[39\] clknet_leaf_111_clk sg13g2_dfrbpq_1
XFILLER_94_217 VPWR VGND sg13g2_fill_2
XFILLER_67_409 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_674 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nand2b_1_B data_pvalid_sg13g2_nand2b_1_B_Y net423 VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[9\]
+ sg13g2_nand2b_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ VPWR VGND sg13g2_and4_2
XFILLER_87_291 VPWR VGND sg13g2_fill_2
XFILLER_76_976 VPWR VGND sg13g2_decap_8
XFILLER_75_464 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2481 i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X
+ net2532 VPWR VGND sg13g2_a22oi_1
XFILLER_36_807 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ net2923 net3034 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A
+ VPWR VGND i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D
+ sg13g2_nand4_1
XFILLER_75_475 VPWR VGND sg13g2_fill_1
XFILLER_47_166 VPWR VGND sg13g2_fill_2
XFILLER_91_968 VPWR VGND sg13g2_decap_8
XFILLER_90_445 VPWR VGND sg13g2_decap_8
XFILLER_35_339 VPWR VGND sg13g2_fill_1
XFILLER_90_489 VPWR VGND sg13g2_decap_8
XFILLER_93_7 VPWR VGND sg13g2_decap_8
XFILLER_43_372 VPWR VGND sg13g2_fill_1
XFILLER_16_597 VPWR VGND sg13g2_decap_8
XFILLER_31_545 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ net2488 i_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D i_snitch.gpr_waddr\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[487\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[487\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2457 net2284 net2367 net1314 VPWR VGND sg13g2_a22oi_1
XFILLER_12_770 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[230\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2287
+ net2437 VPWR VGND sg13g2_nand2_1
XFILLER_7_273 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[382\] clknet_leaf_86_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q
+ net3228 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[171\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[171\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net897 net2679 net2775 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2
+ VGND net2498 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_79_770 VPWR VGND sg13g2_decap_4
Xi_req_register.data_o\[43\]_sg13g2_o21ai_1_Y i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.data_o\[43\] VGND net3166 i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_79_781 VPWR VGND sg13g2_fill_2
XFILLER_67_943 VPWR VGND sg13g2_fill_1
XFILLER_66_420 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2474 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1
+ net86 i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_82_902 VPWR VGND sg13g2_decap_8
XFILLER_15_0 VPWR VGND sg13g2_fill_2
XFILLER_93_250 VPWR VGND sg13g2_fill_2
XFILLER_53_114 VPWR VGND sg13g2_decap_8
XFILLER_26_306 VPWR VGND sg13g2_decap_4
XFILLER_82_979 VPWR VGND sg13g2_decap_8
XFILLER_53_125 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[378\]_sg13g2_o21ai_1_A1 net2968 VPWR i_snitch.i_snitch_regfile.mem\[378\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[378\] net2800 sg13g2_o21ai_1
XFILLER_35_840 VPWR VGND sg13g2_fill_1
Xi_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1 VPWR VGND i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1 net2637 i_req_arb.data_i\[42\] i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y
+ net2721 sg13g2_a221oi_1
XFILLER_50_843 VPWR VGND sg13g2_fill_1
XFILLER_50_832 VPWR VGND sg13g2_decap_8
XFILLER_22_534 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y
+ VGND VPWR net2604 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[201\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[201\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q net3265 VGND VPWR i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[59\] clknet_leaf_113_clk sg13g2_dfrbpq_1
Xhold730 i_snitch.i_snitch_regfile.mem\[460\] VPWR VGND net762 sg13g2_dlygate4sd3_1
XFILLER_104_823 VPWR VGND sg13g2_decap_8
Xhold741 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net773 sg13g2_dlygate4sd3_1
Xhold752 i_snitch.i_snitch_regfile.mem\[503\] VPWR VGND net784 sg13g2_dlygate4sd3_1
Xhold763 i_snitch.i_snitch_regfile.mem\[361\] VPWR VGND net795 sg13g2_dlygate4sd3_1
Xfanout2909 net2910 net2909 VPWR VGND sg13g2_buf_8
XFILLER_103_322 VPWR VGND sg13g2_decap_8
Xhold774 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] VPWR
+ VGND net806 sg13g2_dlygate4sd3_1
Xhold785 i_snitch.i_snitch_regfile.mem\[107\] VPWR VGND net817 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
Xhold796 i_snitch.i_snitch_regfile.mem\[146\] VPWR VGND net828 sg13g2_dlygate4sd3_1
XFILLER_77_718 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1
+ i_req_arb.data_i\[40\] i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_103_399 VPWR VGND sg13g2_decap_8
XFILLER_57_420 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_85_751 VPWR VGND sg13g2_fill_1
XFILLER_58_965 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[6\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]
+ net118 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X
+ VPWR VGND sg13g2_mux2_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 net42 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_and2_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y
+ net2815 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X
+ net3082 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1
+ VPWR VGND sg13g2_and2_1
XFILLER_60_629 VPWR VGND sg13g2_decap_4
XFILLER_38_1023 VPWR VGND sg13g2_decap_4
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net693 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2327 net2892 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_dfrbpq_1_Q_D net2908
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[191\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[191\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2343 net840 net2645 net2773 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[222\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_40_331 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2739 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_X
+ net3095 net2929 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[365\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2291
+ net2470 VPWR VGND sg13g2_nand2_1
XFILLER_84_1010 VPWR VGND sg13g2_decap_8
XFILLER_106_182 VPWR VGND sg13g2_decap_8
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_972 VPWR VGND sg13g2_decap_8
XFILLER_96_63 VPWR VGND sg13g2_decap_8
XFILLER_67_239 VPWR VGND sg13g2_fill_1
XFILLER_67_228 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2740
+ net2669 VPWR VGND sg13g2_nand2_1
XFILLER_0_482 VPWR VGND sg13g2_fill_2
XFILLER_49_965 VPWR VGND sg13g2_fill_1
XFILLER_49_954 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[326\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[326\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2403 net786 net2899 net2796 VPWR VGND sg13g2_a22oi_1
XFILLER_49_987 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_X
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 VPWR VGND
+ sg13g2_nor2_1
XFILLER_63_434 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q net3297 VGND VPWR i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[79\] clknet_leaf_63_clk sg13g2_dfrbpq_1
XFILLER_35_136 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[500\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2845
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[40\]
+ net2826 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y net2821 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[221\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[221\] clknet_leaf_96_clk sg13g2_dfrbpq_1
XFILLER_91_1003 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B
+ i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[2\] net960 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y net110 i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2937 sg13g2_a21oi_1
XFILLER_32_876 VPWR VGND sg13g2_decap_4
XFILLER_105_609 VPWR VGND sg13g2_fill_1
XFILLER_104_119 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[169\]_sg13g2_dfrbpq_1_Q_D VGND net2300 net2340
+ sg13g2_o21ai_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_832 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ net2553 VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B
+ VGND net2715 i_snitch.i_snitch_regfile.mem\[147\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ sg13g2_o21ai_1
Xrsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ net1350 VGND sg13g2_inv_1
XFILLER_58_206 VPWR VGND sg13g2_decap_4
XFILLER_101_826 VPWR VGND sg13g2_decap_8
XFILLER_100_303 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2762 net2307
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1 net2519 sg13g2_a221oi_1
XFILLER_39_420 VPWR VGND sg13g2_fill_1
Xrebuffer11 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y
+ net43 VPWR VGND sg13g2_buf_1
XFILLER_27_626 VPWR VGND sg13g2_fill_2
XFILLER_39_486 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1
+ net557 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xrebuffer33 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y
+ net65 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2708 i_snitch.i_snitch_regfile.mem\[114\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xrebuffer22 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net54 VPWR VGND sg13g2_buf_1
Xrebuffer55 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y
+ net87 VPWR VGND sg13g2_buf_1
XFILLER_82_732 VPWR VGND sg13g2_decap_8
Xrebuffer44 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y
+ net76 VPWR VGND sg13g2_buf_1
XFILLER_66_283 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2413
+ sg13g2_o21ai_1
XFILLER_27_648 VPWR VGND sg13g2_fill_2
Xrebuffer77 net3143 net109 VPWR VGND sg13g2_buf_1
Xrebuffer88 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X
+ net120 VPWR VGND sg13g2_buf_1
Xrebuffer66 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C
+ net98 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1 net2831
+ VPWR i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_dfrbpq_1_Q_D VGND net2276 net2385
+ sg13g2_o21ai_1
XFILLER_23_843 VPWR VGND sg13g2_decap_8
XFILLER_23_898 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1107 net2497 net1269 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[118\]
+ net2806 i_snitch.i_snitch_regfile.mem\[118\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_a22oi_1_B2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2399
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_a22oi_1_B2_Y
+ net2401 net703 net2472 net2255 VPWR VGND sg13g2_a22oi_1
Xfanout2706 net2707 net2706 VPWR VGND sg13g2_buf_8
Xfanout2717 net2718 net2717 VPWR VGND sg13g2_buf_8
Xhold560 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net592 sg13g2_dlygate4sd3_1
Xhold571 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\] VPWR
+ VGND net603 sg13g2_dlygate4sd3_1
XFILLER_2_747 VPWR VGND sg13g2_decap_8
XFILLER_89_364 VPWR VGND sg13g2_fill_1
Xhold582 shift_reg_q\[27\] VPWR VGND net614 sg13g2_dlygate4sd3_1
Xhold593 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\] VPWR
+ VGND net625 sg13g2_dlygate4sd3_1
Xfanout2728 net2729 net2728 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[99\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[99\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[99\] clknet_leaf_100_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nor3_1_A net1219 net2782 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xfanout2739 net2740 net2739 VPWR VGND sg13g2_buf_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[241\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[241\] clknet_leaf_82_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[60\]
+ net2826 i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a21oi_1_A1_Y net2821 sg13g2_a21oi_1
XFILLER_106_84 VPWR VGND sg13g2_decap_8
XFILLER_103_196 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y VPWR VGND net2761 net2310
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2520 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 sg13g2_a221oi_1
XFILLER_58_795 VPWR VGND sg13g2_decap_4
XFILLER_46_924 VPWR VGND sg13g2_decap_8
Xhold1260 i_snitch.i_snitch_regfile.mem\[307\] VPWR VGND net1292 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2415 sg13g2_a21oi_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ net2759 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 VPWR VGND sg13g2_nand2_1
XFILLER_72_220 VPWR VGND sg13g2_decap_8
Xhold1271 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\] VPWR
+ VGND net1303 sg13g2_dlygate4sd3_1
XFILLER_46_957 VPWR VGND sg13g2_decap_4
XFILLER_45_445 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold1293 i_snitch.i_snitch_regfile.mem\[499\] VPWR VGND net1325 sg13g2_dlygate4sd3_1
Xhold1282 i_snitch.i_snitch_regfile.mem\[487\] VPWR VGND net1314 sg13g2_dlygate4sd3_1
XFILLER_73_765 VPWR VGND sg13g2_decap_8
XFILLER_60_415 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[347\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_26_670 VPWR VGND sg13g2_decap_8
XFILLER_32_106 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[5\]_sg13g2_dfrbpq_1_Q net3240 VGND VPWR rsp_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[5\] clknet_leaf_37_clk sg13g2_dfrbpq_2
Xheichips25_snitch_wrapper_26 VPWR VGND uio_oe[6] sg13g2_tiehi
Xi_snitch.i_snitch_regfile.mem\[323\]_sg13g2_nor3_1_A net1311 net2795 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[323\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2571 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ net2539 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y net2846 i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_40_172 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\] net635 net2623
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_Y i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1
+ net2506 i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor3_1_A_C VPWR VGND sg13g2_nor2_2
XFILLER_96_802 VPWR VGND sg13g2_decap_8
XFILLER_68_548 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_nand3b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\] i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[0\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_nand3b_1_B_Y
+ VPWR VGND net3178 sg13g2_nand3b_1
XFILLER_83_518 VPWR VGND sg13g2_decap_8
XFILLER_76_570 VPWR VGND sg13g2_decap_4
XFILLER_48_261 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_dfrbpq_1_Q
+ net3195 VGND VPWR net624 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_36_423 VPWR VGND sg13g2_fill_2
XFILLER_37_968 VPWR VGND sg13g2_fill_2
XFILLER_91_562 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[244\]_sg13g2_dfrbpq_1_Q_D VGND net2260 net2329
+ sg13g2_o21ai_1
XFILLER_36_478 VPWR VGND sg13g2_decap_4
XFILLER_91_584 VPWR VGND sg13g2_fill_2
XFILLER_63_286 VPWR VGND sg13g2_fill_2
XFILLER_52_949 VPWR VGND sg13g2_fill_2
XFILLER_51_448 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net1194 net2687 net2881 VPWR VGND sg13g2_a22oi_1
XFILLER_32_695 VPWR VGND sg13g2_decap_8
XFILLER_9_880 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A
+ sg13g2_or2_1
XFILLER_11_28 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[80\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[80\]
+ net2844 i_snitch.i_snitch_regfile.mem\[80\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q net3218 VGND VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[261\] clknet_leaf_110_clk sg13g2_dfrbpq_1
XFILLER_105_406 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2585 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2377
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_A
+ net2703 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[367\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[367\]
+ net3135 i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_a21oi_1_A1_Y net2944 sg13g2_a21oi_1
XFILLER_101_601 VPWR VGND sg13g2_decap_4
XFILLER_99_695 VPWR VGND sg13g2_fill_1
XFILLER_59_526 VPWR VGND sg13g2_fill_1
XFILLER_101_656 VPWR VGND sg13g2_fill_1
XFILLER_100_133 VPWR VGND sg13g2_decap_8
XFILLER_100_177 VPWR VGND sg13g2_decap_8
XFILLER_86_378 VPWR VGND sg13g2_fill_1
XFILLER_86_367 VPWR VGND sg13g2_fill_2
XFILLER_74_529 VPWR VGND sg13g2_fill_1
XFILLER_28_968 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[372\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[340\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2828
+ sg13g2_a221oi_1
XFILLER_55_765 VPWR VGND sg13g2_decap_4
XFILLER_82_584 VPWR VGND sg13g2_fill_2
XFILLER_74_1020 VPWR VGND sg13g2_decap_8
XFILLER_70_746 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ net2518 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ net2755 VPWR VGND sg13g2_a22oi_1
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_42_426 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[268\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[364\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2846
+ sg13g2_a221oi_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y
+ VPWR VGND sg13g2_and3_2
XFILLER_10_367 VPWR VGND sg13g2_decap_4
XFILLER_10_345 VPWR VGND sg13g2_decap_8
Xfanout3204 net3205 net3204 VPWR VGND sg13g2_buf_2
Xfanout3237 net3239 net3237 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]_sg13g2_dfrbpq_1_Q
+ net3203 VGND VPWR net433 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[36\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_1
Xfanout3215 net3216 net3215 VPWR VGND sg13g2_buf_8
XFILLER_2_511 VPWR VGND sg13g2_decap_8
Xfanout3226 net3330 net3226 VPWR VGND sg13g2_buf_8
XFILLER_105_973 VPWR VGND sg13g2_decap_8
Xfanout3248 net3249 net3248 VPWR VGND sg13g2_buf_8
Xfanout2525 net2529 net2525 VPWR VGND sg13g2_buf_8
Xfanout2536 net2536 net2537 VPWR VGND sg13g2_buf_16
Xfanout3259 net3261 net3259 VPWR VGND sg13g2_buf_8
Xfanout2514 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_Y
+ net2514 VPWR VGND sg13g2_buf_8
Xfanout2503 net2505 net2503 VPWR VGND sg13g2_buf_8
Xfanout2558 net2559 net2558 VPWR VGND sg13g2_buf_1
Xfanout2547 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y
+ net2547 VPWR VGND sg13g2_buf_8
Xfanout2569 net2570 net2569 VPWR VGND sg13g2_buf_8
XFILLER_2_577 VPWR VGND sg13g2_fill_1
XFILLER_77_367 VPWR VGND sg13g2_decap_8
XFILLER_93_42 VPWR VGND sg13g2_decap_8
XFILLER_92_326 VPWR VGND sg13g2_decap_4
XFILLER_45_220 VPWR VGND sg13g2_fill_1
Xhold1090 i_snitch.wake_up_q\[0\] VPWR VGND net1122 sg13g2_dlygate4sd3_1
XFILLER_73_573 VPWR VGND sg13g2_fill_1
XFILLER_61_735 VPWR VGND sg13g2_decap_8
XFILLER_45_264 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q net3216 VGND VPWR i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[281\] clknet_leaf_115_clk sg13g2_dfrbpq_1
XFILLER_60_289 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2628 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1
+ net2755 VPWR VGND sg13g2_a22oi_1
Xrebuffer2 net33 net34 VPWR VGND sg13g2_buf_2
XFILLER_61_5 VPWR VGND sg13g2_fill_1
XFILLER_6_872 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[416\] clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_68_323 VPWR VGND sg13g2_fill_1
XFILLER_56_529 VPWR VGND sg13g2_fill_2
XFILLER_56_518 VPWR VGND sg13g2_fill_1
XFILLER_3_84 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[205\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[205\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2338 net1041 net2690 net2792 VPWR VGND sg13g2_a22oi_1
XFILLER_97_1020 VPWR VGND sg13g2_decap_8
XFILLER_84_849 VPWR VGND sg13g2_decap_8
XFILLER_92_871 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_nor2b_1_B_N
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_nor2b_1
XFILLER_51_212 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q net3223 VGND VPWR i_snitch.i_snitch_regfile.mem\[100\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[100\] clknet_leaf_106_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A_Y net2952 i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2944 sg13g2_a21oi_1
XFILLER_33_960 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2631 VPWR i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1
+ net2751 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_mux2_1_A1_1_X
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_dfrbpq_1_Q net3252 VGND VPWR i_snitch.i_snitch_lsu.handshake_pending_d
+ i_snitch.i_snitch_lsu.handshake_pending_q clknet_leaf_21_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ sg13g2_nand2b_2
XFILLER_106_759 VPWR VGND sg13g2_decap_8
XFILLER_105_203 VPWR VGND sg13g2_decap_8
XFILLER_99_470 VPWR VGND sg13g2_fill_1
XFILLER_87_610 VPWR VGND sg13g2_fill_2
XFILLER_59_301 VPWR VGND sg13g2_fill_2
XFILLER_102_954 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] net603 net2621
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_101_475 VPWR VGND sg13g2_fill_2
XFILLER_59_367 VPWR VGND sg13g2_fill_1
XFILLER_59_356 VPWR VGND sg13g2_decap_8
XFILLER_75_849 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2
+ VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A i_snitch.inst_addr_o\[15\]
+ net2527 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A net2535
+ net3071 i_snitch.inst_addr_o\[1\] VPWR VGND sg13g2_and3_1
Xshift_reg_q\[7\]_sg13g2_dfrbpq_1_Q net3195 VGND VPWR net493 shift_reg_q\[7\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_103_63 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2582 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_83_893 VPWR VGND sg13g2_decap_8
XFILLER_82_370 VPWR VGND sg13g2_fill_1
XFILLER_70_521 VPWR VGND sg13g2_decap_8
XFILLER_55_573 VPWR VGND sg13g2_fill_1
XFILLER_42_223 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0 net3138 i_snitch.i_snitch_regfile.mem\[150\]
+ i_snitch.i_snitch_regfile.mem\[182\] i_snitch.i_snitch_regfile.mem\[214\] i_snitch.i_snitch_regfile.mem\[246\]
+ net3111 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y
+ net2533 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2697 i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2
+ net2541 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[297\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[297\] net2811 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[436\] clknet_leaf_59_clk sg13g2_dfrbpq_1
XFILLER_7_658 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B
+ VPWR VGND i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N
+ sg13g2_nand3b_1
XFILLER_12_71 VPWR VGND sg13g2_fill_1
Xfanout3012 net3015 net3012 VPWR VGND sg13g2_buf_8
Xfanout3001 net3003 net3001 VPWR VGND sg13g2_buf_8
Xfanout3034 net3037 net3034 VPWR VGND sg13g2_buf_8
Xfanout2311 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B_X
+ net2311 VPWR VGND sg13g2_buf_8
Xfanout3023 net3024 net3023 VPWR VGND sg13g2_buf_8
Xfanout2300 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2300 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_X
+ net3096 net2931 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_3_864 VPWR VGND sg13g2_decap_8
Xfanout3045 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X net3045 VPWR VGND sg13g2_buf_8
XFILLER_105_770 VPWR VGND sg13g2_decap_8
XFILLER_97_429 VPWR VGND sg13g2_decap_4
Xfanout3078 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1_1_X
+ net3078 VPWR VGND sg13g2_buf_8
Xfanout3067 rsp_data_ready net3067 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q net3324 VGND VPWR i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[120\] clknet_leaf_58_clk sg13g2_dfrbpq_1
Xfanout3089 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_mux2_1_A1_X
+ net3089 VPWR VGND sg13g2_buf_8
Xfanout3056 state_sg13g2_inv_1_A_Y net3056 VPWR VGND sg13g2_buf_8
Xfanout2344 net2346 net2344 VPWR VGND sg13g2_buf_8
Xfanout2333 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2333 VPWR VGND sg13g2_buf_8
Xfanout2322 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2322 VPWR VGND sg13g2_buf_8
XFILLER_104_280 VPWR VGND sg13g2_decap_8
Xfanout2366 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2366 VPWR VGND sg13g2_buf_8
Xfanout2377 net2378 net2377 VPWR VGND sg13g2_buf_8
Xfanout2355 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2355 VPWR VGND sg13g2_buf_8
XFILLER_66_816 VPWR VGND sg13g2_decap_8
Xfanout2399 net2400 net2399 VPWR VGND sg13g2_buf_8
Xfanout2388 i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2388 VPWR VGND sg13g2_buf_8
XFILLER_93_624 VPWR VGND sg13g2_fill_2
XFILLER_19_732 VPWR VGND sg13g2_fill_2
XFILLER_92_167 VPWR VGND sg13g2_fill_1
XFILLER_65_359 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1 i_snitch.inst_addr_o\[19\] VPWR VGND sg13g2_nand2_2
XFILLER_61_554 VPWR VGND sg13g2_fill_1
XFILLER_22_908 VPWR VGND sg13g2_decap_8
XFILLER_33_267 VPWR VGND sg13g2_fill_2
XFILLER_61_598 VPWR VGND sg13g2_decap_4
XFILLER_88_1008 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[17\]_sg13g2_dfrbpq_1_Q net3231 VGND VPWR rsp_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[17\] clknet_leaf_35_clk sg13g2_dfrbpq_2
XFILLER_6_680 VPWR VGND sg13g2_fill_1
XFILLER_88_407 VPWR VGND sg13g2_decap_8
XFILLER_102_217 VPWR VGND sg13g2_decap_8
XFILLER_97_985 VPWR VGND sg13g2_decap_8
XFILLER_96_473 VPWR VGND sg13g2_fill_2
XFILLER_96_451 VPWR VGND sg13g2_fill_2
XFILLER_84_602 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ net2550 VPWR i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ VGND i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ net2715 sg13g2_o21ai_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1
+ VPWR VGND sg13g2_nand2_1
XFILLER_84_624 VPWR VGND sg13g2_decap_8
XFILLER_25_724 VPWR VGND sg13g2_decap_8
XFILLER_80_830 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q net3280 VGND VPWR i_snitch.i_snitch_regfile.mem\[456\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[456\] clknet_leaf_74_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[322\] net2947 VPWR VGND sg13g2_nand2_1
XFILLER_80_896 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ net2993 net2725 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[245\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[245\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2330 net1095 net2438 net2268 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2557 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q net3310 VGND VPWR i_snitch.i_snitch_regfile.mem\[140\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[140\] clknet_leaf_68_clk sg13g2_dfrbpq_1
XFILLER_20_462 VPWR VGND sg13g2_fill_1
XFILLER_20_473 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ net2628 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ net2756 VPWR VGND sg13g2_a22oi_1
XFILLER_4_617 VPWR VGND sg13g2_fill_2
XFILLER_106_523 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_88_952 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[403\] net3026 VPWR VGND sg13g2_nand2_1
XFILLER_0_856 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VGND sg13g2_inv_1
XFILLER_87_473 VPWR VGND sg13g2_fill_2
XFILLER_75_613 VPWR VGND sg13g2_fill_2
XFILLER_47_304 VPWR VGND sg13g2_decap_8
XFILLER_87_484 VPWR VGND sg13g2_fill_2
XFILLER_75_635 VPWR VGND sg13g2_fill_2
XFILLER_101_294 VPWR VGND sg13g2_decap_8
XFILLER_74_156 VPWR VGND sg13g2_fill_2
XFILLER_47_359 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1
+ VGND VPWR net3078 net2850 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ sg13g2_a21oi_1
XFILLER_74_55 VPWR VGND sg13g2_fill_2
XFILLER_90_21 VPWR VGND sg13g2_decap_8
XFILLER_71_874 VPWR VGND sg13g2_decap_4
XFILLER_70_351 VPWR VGND sg13g2_decap_8
XFILLER_16_779 VPWR VGND sg13g2_decap_4
XFILLER_24_790 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2
+ net41 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_a21o_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_7_433 VPWR VGND sg13g2_decap_8
XFILLER_7_411 VPWR VGND sg13g2_fill_2
XFILLER_23_81 VPWR VGND sg13g2_decap_4
XFILLER_7_455 VPWR VGND sg13g2_fill_2
XFILLER_99_63 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND net2703 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ net2545 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2415 i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_66_602 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q net3267 VGND VPWR i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[476\] clknet_leaf_96_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_a22oi_1_B2_Y
+ net2327 net644 net2685 net2892 VPWR VGND sg13g2_a22oi_1
XFILLER_94_966 VPWR VGND sg13g2_decap_8
XFILLER_94_1001 VPWR VGND sg13g2_decap_8
XFILLER_65_189 VPWR VGND sg13g2_decap_8
XFILLER_46_370 VPWR VGND sg13g2_fill_1
XFILLER_34_510 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q net3256 VGND VPWR i_snitch.i_snitch_regfile.mem\[160\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[160\] clknet_leaf_49_clk sg13g2_dfrbpq_1
XFILLER_0_63 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[107\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ net2531 i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[342\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0 net3126 i_snitch.i_snitch_regfile.mem\[157\]
+ i_snitch.i_snitch_regfile.mem\[189\] i_snitch.i_snitch_regfile.mem\[221\] i_snitch.i_snitch_regfile.mem\[253\]
+ net3106 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 net2627 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A_Y
+ net2758 VPWR VGND sg13g2_a22oi_1
Xhold901 i_snitch.i_snitch_regfile.mem\[447\] VPWR VGND net933 sg13g2_dlygate4sd3_1
Xhold912 i_snitch.i_snitch_regfile.mem\[278\] VPWR VGND net944 sg13g2_dlygate4sd3_1
Xdata_pdata\[18\]_sg13g2_dfrbpq_1_Q net3201 VGND VPWR net750 data_pdata\[18\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
Xhold923 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net955 sg13g2_dlygate4sd3_1
Xhold934 data_pdata\[15\] VPWR VGND net966 sg13g2_dlygate4sd3_1
Xhold945 i_snitch.i_snitch_regfile.mem\[79\] VPWR VGND net977 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net463 net2350 VPWR VGND sg13g2_nand2_1
XFILLER_103_504 VPWR VGND sg13g2_decap_4
Xhold967 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net999 sg13g2_dlygate4sd3_1
XFILLER_89_727 VPWR VGND sg13g2_fill_2
Xhold956 i_snitch.i_snitch_regfile.mem\[371\] VPWR VGND net988 sg13g2_dlygate4sd3_1
Xhold989 i_snitch.i_snitch_regfile.mem\[378\] VPWR VGND net1021 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[208\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold978 i_snitch.i_snitch_regfile.mem\[82\] VPWR VGND net1010 sg13g2_dlygate4sd3_1
XFILLER_103_537 VPWR VGND sg13g2_fill_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0_X
+ net2939 net2929 i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_96_270 VPWR VGND sg13g2_fill_2
XFILLER_85_955 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_48 VPWR VGND sg13g2_fill_1
XFILLER_29_326 VPWR VGND sg13g2_fill_1
XFILLER_38_871 VPWR VGND sg13g2_fill_2
XFILLER_38_893 VPWR VGND sg13g2_fill_2
XFILLER_52_340 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_100_42 VPWR VGND sg13g2_decap_8
XFILLER_21_771 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q net3290 VGND VPWR i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[496\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_20_281 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2324 net884 net2434 net2251 VPWR VGND sg13g2_a22oi_1
XFILLER_106_364 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[35\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y
+ net2479 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2530 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[180\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[180\] clknet_leaf_56_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[178\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_653 VPWR VGND sg13g2_decap_8
XFILLER_91_947 VPWR VGND sg13g2_decap_8
XFILLER_29_860 VPWR VGND sg13g2_decap_4
Xrsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1107 net3065 rsp_data_q\[27\] VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y
+ net1393 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_16_521 VPWR VGND sg13g2_decap_8
XFILLER_18_92 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2
+ VGND net2712 i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_565 VPWR VGND sg13g2_fill_1
XFILLER_71_682 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[472\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[329\] net2949 VPWR VGND sg13g2_nand2_1
XFILLER_86_7 VPWR VGND sg13g2_fill_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q net3235 VGND VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D
+ i_req_arb.gen_arbiter.rr_q clknet_leaf_22_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0 net3021 i_snitch.i_snitch_regfile.mem\[395\]
+ i_snitch.i_snitch_regfile.mem\[427\] i_snitch.i_snitch_regfile.mem\[459\] i_snitch.i_snitch_regfile.mem\[491\]
+ net2992 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
XFILLER_8_742 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q net3214 VGND VPWR i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[315\] clknet_leaf_117_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[104\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2410 net849 net2643 net2869 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2443 net2772 i_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q_D net2909
+ sg13g2_a221oi_1
XFILLER_98_524 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2
+ net2614 i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[22\]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_a21o_1
XFILLER_86_708 VPWR VGND sg13g2_fill_2
XFILLER_38_112 VPWR VGND sg13g2_fill_1
XFILLER_94_741 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_inv_1_A
+ VPWR data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y
+ VGND sg13g2_inv_1
XFILLER_93_262 VPWR VGND sg13g2_fill_1
Xdata_pdata\[23\]_sg13g2_mux2_1_A1 rsp_data_q\[23\] net721 net3050 data_pdata\[23\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_82_958 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net73 net2851 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A_Y
+ sg13g2_a21oi_1
XFILLER_81_446 VPWR VGND sg13g2_fill_2
XFILLER_53_148 VPWR VGND sg13g2_fill_1
XFILLER_81_479 VPWR VGND sg13g2_decap_8
XFILLER_81_468 VPWR VGND sg13g2_fill_2
XFILLER_53_159 VPWR VGND sg13g2_decap_8
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_90_980 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_nand2_1_A_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[41\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.data_o\[41\]_sg13g2_o21ai_1_Y_A2 net2616 sg13g2_o21ai_1
Xhold720 i_snitch.i_snitch_regfile.mem\[136\] VPWR VGND net752 sg13g2_dlygate4sd3_1
XFILLER_104_802 VPWR VGND sg13g2_decap_8
Xhold731 i_req_arb.gen_arbiter.rr_q VPWR VGND net763 sg13g2_dlygate4sd3_1
Xhold764 i_snitch.i_snitch_regfile.mem\[440\] VPWR VGND net796 sg13g2_dlygate4sd3_1
Xhold753 i_snitch.i_snitch_regfile.mem\[276\] VPWR VGND net785 sg13g2_dlygate4sd3_1
XFILLER_2_929 VPWR VGND sg13g2_decap_8
Xhold742 i_snitch.i_snitch_regfile.mem\[465\] VPWR VGND net774 sg13g2_dlygate4sd3_1
XFILLER_103_301 VPWR VGND sg13g2_decap_8
XFILLER_89_557 VPWR VGND sg13g2_fill_2
XFILLER_89_546 VPWR VGND sg13g2_decap_8
Xhold775 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net807 sg13g2_dlygate4sd3_1
Xhold797 i_snitch.i_snitch_regfile.mem\[431\] VPWR VGND net829 sg13g2_dlygate4sd3_1
Xhold786 data_pdata\[26\] VPWR VGND net818 sg13g2_dlygate4sd3_1
XFILLER_104_879 VPWR VGND sg13g2_decap_8
XFILLER_89_579 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_103_378 VPWR VGND sg13g2_decap_8
XFILLER_58_944 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[217\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2788
+ net2661 VPWR VGND sg13g2_nand2_1
XFILLER_29_112 VPWR VGND sg13g2_fill_2
XFILLER_57_454 VPWR VGND sg13g2_fill_2
XFILLER_57_432 VPWR VGND sg13g2_fill_2
XFILLER_85_774 VPWR VGND sg13g2_decap_4
XFILLER_84_273 VPWR VGND sg13g2_fill_1
XFILLER_73_947 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[335\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[335\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2838 i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q
+ net3252 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[502\]_sg13g2_o21ai_1_A1 net2965 VPWR i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[502\] net2806 sg13g2_o21ai_1
XFILLER_81_991 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[124\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[124\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2449 net2247 net2409 net1201 VPWR VGND sg13g2_a22oi_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B i_snitch.gpr_waddr\[7\]_sg13g2_nor2_1_A_Y
+ data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X
+ VPWR VGND sg13g2_and2_1
XFILLER_41_811 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
XFILLER_9_506 VPWR VGND sg13g2_decap_8
XFILLER_9_517 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[253\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1
+ net2684 i_snitch.i_snitch_regfile.mem\[154\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_71_78 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nor2b_1
Xshift_reg_q\[23\]_sg13g2_a22oi_1_A1 shift_reg_q\[23\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_mux2_1_A1_1_X
+ net3056 net3046 shift_reg_q\[23\] VPWR VGND sg13g2_a22oi_1
XFILLER_5_789 VPWR VGND sg13g2_fill_2
XFILLER_106_161 VPWR VGND sg13g2_decap_8
XFILLER_96_42 VPWR VGND sg13g2_decap_8
XFILLER_68_719 VPWR VGND sg13g2_fill_2
XFILLER_68_708 VPWR VGND sg13g2_decap_8
XFILLER_1_951 VPWR VGND sg13g2_decap_8
XFILLER_0_461 VPWR VGND sg13g2_decap_8
XFILLER_64_903 VPWR VGND sg13g2_fill_2
XFILLER_49_977 VPWR VGND sg13g2_fill_1
XFILLER_48_443 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2543 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2889
+ net2667 VPWR VGND sg13g2_nand2_1
XFILLER_29_91 VPWR VGND sg13g2_fill_1
XFILLER_91_744 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[457\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2378
+ sg13g2_o21ai_1
XFILLER_17_841 VPWR VGND sg13g2_decap_8
XFILLER_63_479 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[270\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2725 i_snitch.inst_addr_o\[14\] sg13g2_a21oi_2
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net2928 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_C1 net70 i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1
+ sg13g2_a21oi_2
XFILLER_71_490 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_70_clk clknet_5_25__leaf_clk clknet_leaf_70_clk VPWR VGND sg13g2_buf_8
XFILLER_99_811 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2431
+ net2291 VPWR VGND sg13g2_nand2_1
XFILLER_101_805 VPWR VGND sg13g2_decap_8
XFILLER_99_888 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ net2587 i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[355\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[355\] clknet_leaf_108_clk sg13g2_dfrbpq_1
XFILLER_98_398 VPWR VGND sg13g2_fill_2
XFILLER_100_359 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net1047 net2446 net2262 VPWR VGND sg13g2_a22oi_1
XFILLER_94_560 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y i_snitch.pc_d\[16\] i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2 net2308 i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
Xrebuffer12 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y
+ net44 VPWR VGND sg13g2_buf_2
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2347
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_and2_1_X
+ net2923 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2
+ VPWR VGND sg13g2_and2_1
Xrebuffer23 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ net55 VPWR VGND sg13g2_buf_2
Xrebuffer45 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A
+ net77 VPWR VGND sg13g2_buf_1
Xrebuffer34 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ net66 VPWR VGND sg13g2_buf_1
XFILLER_66_295 VPWR VGND sg13g2_fill_2
XFILLER_55_947 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2669 VPWR VGND sg13g2_nand2_1
Xrebuffer56 net2563 net88 VPWR VGND sg13g2_buf_1
Xrebuffer67 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B
+ net99 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2638 i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
Xrebuffer78 net2921 net110 VPWR VGND sg13g2_buf_1
Xrebuffer89 net3181 net121 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_61_clk clknet_5_29__leaf_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ net2924 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_a22oi_1
XFILLER_68_1028 VPWR VGND sg13g2_fill_1
XFILLER_68_1017 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_B1
+ net695 net2767 VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[509\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2858
+ net2653 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B
+ net2640 i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_2
XFILLER_104_610 VPWR VGND sg13g2_fill_1
Xfanout2707 net2708 net2707 VPWR VGND sg13g2_buf_8
XFILLER_89_332 VPWR VGND sg13g2_decap_4
Xfanout2718 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N_Y
+ net2718 VPWR VGND sg13g2_buf_8
Xi_snitch.inst_addr_o\[15\]_sg13g2_dfrbpq_1_Q net3327 VGND VPWR i_snitch.pc_d\[15\]
+ i_snitch.inst_addr_o\[15\] clknet_leaf_58_clk sg13g2_dfrbpq_2
Xhold572 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net604 sg13g2_dlygate4sd3_1
Xhold561 i_snitch.sb_q\[3\] VPWR VGND net593 sg13g2_dlygate4sd3_1
Xhold550 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\] VPWR
+ VGND net582 sg13g2_dlygate4sd3_1
XFILLER_2_726 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xhold583 shift_reg_q\[27\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net615 sg13g2_dlygate4sd3_1
Xhold594 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[25\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net626 sg13g2_dlygate4sd3_1
Xfanout2729 net2730 net2729 VPWR VGND sg13g2_buf_8
XFILLER_106_63 VPWR VGND sg13g2_decap_8
XFILLER_103_175 VPWR VGND sg13g2_decap_8
XFILLER_89_398 VPWR VGND sg13g2_decap_8
XFILLER_66_45 VPWR VGND sg13g2_fill_2
XFILLER_58_741 VPWR VGND sg13g2_decap_8
XFILLER_100_882 VPWR VGND sg13g2_decap_8
Xhold1261 rsp_data_q\[29\] VPWR VGND net1293 sg13g2_dlygate4sd3_1
XFILLER_45_402 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[305\]_sg13g2_dfrbpq_1_Q_D VGND net2314 net2288
+ sg13g2_o21ai_1
Xhold1250 i_snitch.i_snitch_regfile.mem\[162\] VPWR VGND net1282 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2
+ VPWR VGND net2544 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ net2699 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ sg13g2_a221oi_1
XFILLER_85_582 VPWR VGND sg13g2_fill_1
XFILLER_73_722 VPWR VGND sg13g2_fill_2
XFILLER_45_435 VPWR VGND sg13g2_fill_1
Xhold1272 i_snitch.i_snitch_regfile.mem\[293\] VPWR VGND net1304 sg13g2_dlygate4sd3_1
Xhold1294 i_snitch.i_snitch_regfile.mem\[34\] VPWR VGND net1326 sg13g2_dlygate4sd3_1
Xhold1283 i_snitch.i_snitch_regfile.mem\[420\] VPWR VGND net1315 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y
+ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_52_clk clknet_5_26__leaf_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
Xheichips25_snitch_wrapper_27 VPWR VGND uio_oe[5] sg13g2_tiehi
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]_sg13g2_dfrbpq_1_Q
+ net3241 VGND VPWR net1019 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[4\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_A2_sg13g2_nor2_1_Y net3127
+ net3106 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_A2 VPWR VGND sg13g2_nor2_2
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q net3310 VGND VPWR i_snitch.i_snitch_regfile.mem\[375\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[375\] clknet_leaf_69_clk sg13g2_dfrbpq_1
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2
+ VGND VPWR net3167 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A_Y
+ strb_reg_q\[0\]_sg13g2_a22oi_1_A1_B2 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1
+ sg13g2_a21oi_1
XFILLER_5_542 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2564 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[36\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[33\]_sg13g2_nand2_1_A_1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_1_Y
+ sg13g2_o21ai_1
XFILLER_95_302 VPWR VGND sg13g2_fill_1
XFILLER_49_752 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2739
+ i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1
+ net570 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
XFILLER_49_774 VPWR VGND sg13g2_decap_8
XFILLER_52_906 VPWR VGND sg13g2_decap_4
XFILLER_63_298 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_43_clk clknet_5_15__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2418 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1 VPWR
+ VGND net2833 net2639 i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1_Y net2954
+ i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y i_snitch.i_snitch_regfile.mem\[397\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y
+ sg13g2_a221oi_1
XFILLER_31_140 VPWR VGND sg13g2_decap_4
XFILLER_75_0 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2335
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2296 net1306 net2494 net1240 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_86_313 VPWR VGND sg13g2_decap_8
XFILLER_100_112 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VGND net75 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ sg13g2_o21ai_1
XFILLER_101_668 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[194\]_sg13g2_nor3_1_A net1238 net2788 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[194\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_27_435 VPWR VGND sg13g2_fill_2
XFILLER_82_552 VPWR VGND sg13g2_decap_8
XFILLER_54_243 VPWR VGND sg13g2_fill_1
XFILLER_43_917 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q
+ net3190 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q net3316 VGND VPWR i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[395\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2738
+ net2673 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_34_clk clknet_5_11__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[184\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net790 net2665 net2775 VPWR VGND sg13g2_a22oi_1
XFILLER_23_630 VPWR VGND sg13g2_decap_4
XFILLER_35_1016 VPWR VGND sg13g2_decap_8
XFILLER_35_1027 VPWR VGND sg13g2_fill_2
XFILLER_50_471 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[184\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2341
+ sg13g2_o21ai_1
XFILLER_10_379 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2360 net861 net2904 net2767 VPWR VGND sg13g2_a22oi_1
Xfanout3238 net3239 net3238 VPWR VGND sg13g2_buf_8
Xfanout3227 net3229 net3227 VPWR VGND sg13g2_buf_8
Xfanout3216 net3226 net3216 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A_Y net3014 sg13g2_o21ai_1
Xfanout3205 net3226 net3205 VPWR VGND sg13g2_buf_8
XFILLER_105_952 VPWR VGND sg13g2_decap_8
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_or2_1_X
+ VGND VPWR i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ sg13g2_or2_1
Xfanout2526 net2529 net2526 VPWR VGND sg13g2_buf_1
Xfanout2515 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y
+ net2515 VPWR VGND sg13g2_buf_8
Xfanout3249 net3330 net3249 VPWR VGND sg13g2_buf_8
Xfanout2504 net2505 net2504 VPWR VGND sg13g2_buf_1
Xfanout2559 net2560 net2559 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2542 VPWR i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1
+ VGND net2750 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xfanout2548 i_snitch.i_snitch_regfile.mem\[438\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2548 VPWR VGND sg13g2_buf_8
Xfanout2537 net2537 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X
+ VPWR VGND sg13g2_buf_16
Xhold391 data_pvalid VPWR VGND net423 sg13g2_dlygate4sd3_1
XFILLER_2_589 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[319\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[319\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2645 net2780 net2318 net1232 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2749 i_snitch.i_snitch_regfile.mem\[400\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_93_839 VPWR VGND sg13g2_decap_8
XFILLER_93_21 VPWR VGND sg13g2_decap_8
Xi_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1
+ i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 net3072 i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_18_435 VPWR VGND sg13g2_fill_2
XFILLER_19_947 VPWR VGND sg13g2_fill_1
XFILLER_73_552 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q net3322 VGND VPWR i_snitch.i_snitch_regfile.mem\[214\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[214\] clknet_leaf_61_clk sg13g2_dfrbpq_1
Xhold1080 i_snitch.i_snitch_regfile.mem\[492\] VPWR VGND net1112 sg13g2_dlygate4sd3_1
Xhold1091 i_snitch.i_snitch_regfile.mem\[466\] VPWR VGND net1123 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[477\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[477\] VGND sg13g2_inv_1
XFILLER_46_788 VPWR VGND sg13g2_fill_1
XFILLER_33_427 VPWR VGND sg13g2_fill_1
XFILLER_61_769 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_25_clk clknet_5_9__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2363
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3040
+ net2694 VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1_sg13g2_or2_1_X
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\] net3179 sg13g2_or2_1
Xstrb_reg_q\[3\]_sg13g2_a21oi_1_A1 VGND VPWR net459 net3043 strb_reg_q\[3\]_sg13g2_a21oi_1_A1_Y
+ strb_reg_q\[2\]_sg13g2_a21oi_1_A1_B1 sg13g2_a21oi_1
Xrebuffer3 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y
+ net35 VPWR VGND sg13g2_buf_8
XFILLER_47_4 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2858
+ net2675 VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net3176 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[23\]
+ sg13g2_o21ai_1
XFILLER_3_63 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_96_699 VPWR VGND sg13g2_fill_2
XFILLER_68_379 VPWR VGND sg13g2_fill_2
XFILLER_68_368 VPWR VGND sg13g2_fill_2
XFILLER_83_327 VPWR VGND sg13g2_decap_8
XFILLER_77_880 VPWR VGND sg13g2_fill_2
XFILLER_49_571 VPWR VGND sg13g2_decap_4
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
XFILLER_92_850 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[420\]_sg13g2_nor3_1_A net1315 net2861 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[420\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xrsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ net1344 VGND sg13g2_inv_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_mux2_1_A1
+ net706 net559 net2238 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_16_clk clknet_5_7__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_mux2_1_A0_X net3114 net2828 i_snitch.i_snitch_regfile.mem\[52\]
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2362 net880 net2672 net2769 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A
+ net116 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_mux2_1_A1_1_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ VPWR VGND sg13g2_nor2b_2
XFILLER_60_791 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2 net2833
+ VPWR i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a22oi_1_A1_Y
+ sg13g2_o21ai_1
Xdata_pdata\[22\]_sg13g2_nor2b_1_B_N net3162 data_pdata\[22\] data_pdata\[22\]_sg13g2_nor2b_1_B_N_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.i_snitch_regfile.mem\[339\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[339\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net1070 net2472 net2271 VPWR VGND sg13g2_a22oi_1
XFILLER_106_727 VPWR VGND sg13g2_decap_8
XFILLER_105_259 VPWR VGND sg13g2_decap_8
XFILLER_59_313 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[53\]
+ net2825 i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a21oi_1_A1_Y net2821 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q net3278 VGND VPWR i_snitch.i_snitch_regfile.mem\[234\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[234\] clknet_leaf_94_clk sg13g2_dfrbpq_1
XFILLER_102_933 VPWR VGND sg13g2_decap_8
XFILLER_101_432 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C
+ i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_87_633 VPWR VGND sg13g2_decap_8
XFILLER_87_688 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A i_snitch.inst_addr_o\[11\]
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_B_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[98\]_sg13g2_nor2_1_A_B
+ net3016 net2989 VPWR VGND sg13g2_nand2_1
XFILLER_68_891 VPWR VGND sg13g2_fill_2
XFILLER_103_42 VPWR VGND sg13g2_decap_8
XFILLER_28_766 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y
+ VPWR VGND sg13g2_and3_2
XFILLER_83_872 VPWR VGND sg13g2_decap_8
XFILLER_70_500 VPWR VGND sg13g2_fill_2
XFILLER_28_799 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X
+ net39 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_xor2_1
XFILLER_82_393 VPWR VGND sg13g2_fill_1
XFILLER_63_46 VPWR VGND sg13g2_decap_4
XFILLER_55_596 VPWR VGND sg13g2_decap_8
XFILLER_63_68 VPWR VGND sg13g2_fill_2
XFILLER_42_279 VPWR VGND sg13g2_decap_8
XFILLER_11_644 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]
+ net3164 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[333\] VGND sg13g2_inv_1
Xfanout3002 net3003 net3002 VPWR VGND sg13g2_buf_1
Xfanout3013 net3015 net3013 VPWR VGND sg13g2_buf_8
Xfanout3035 net3037 net3035 VPWR VGND sg13g2_buf_2
XFILLER_88_43 VPWR VGND sg13g2_decap_8
Xfanout2301 net2302 net2301 VPWR VGND sg13g2_buf_8
Xfanout3024 net3025 net3024 VPWR VGND sg13g2_buf_8
Xfanout3046 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X net3046 VPWR VGND sg13g2_buf_8
XFILLER_3_843 VPWR VGND sg13g2_decap_8
Xfanout3079 net3080 net3079 VPWR VGND sg13g2_buf_8
Xfanout2312 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ net2312 VPWR VGND sg13g2_buf_8
Xfanout3057 state_sg13g2_inv_1_A_Y net3057 VPWR VGND sg13g2_buf_1
Xfanout2334 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2334 VPWR VGND sg13g2_buf_8
Xfanout2323 net2327 net2323 VPWR VGND sg13g2_buf_8
Xfanout3068 net3069 net3068 VPWR VGND sg13g2_buf_8
XFILLER_78_644 VPWR VGND sg13g2_fill_1
Xfanout2367 net2371 net2367 VPWR VGND sg13g2_buf_8
Xdata_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[14\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[30\]_sg13g2_nand2b_1_B_Y net3154 data_pdata\[22\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[14\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
Xfanout2345 net2346 net2345 VPWR VGND sg13g2_buf_8
Xfanout2378 i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ net2378 VPWR VGND sg13g2_buf_8
Xfanout2356 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2356 VPWR VGND sg13g2_buf_8
XFILLER_78_666 VPWR VGND sg13g2_decap_8
Xfanout2389 net2391 net2389 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[17\] net1042 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[72\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[72\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2354 net900 net2643 net2785 VPWR VGND sg13g2_a22oi_1
XFILLER_74_850 VPWR VGND sg13g2_fill_2
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_19_744 VPWR VGND sg13g2_decap_4
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_73_360 VPWR VGND sg13g2_fill_2
XFILLER_46_585 VPWR VGND sg13g2_fill_2
XFILLER_18_254 VPWR VGND sg13g2_fill_1
XFILLER_37_80 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2696 net2548 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[359\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net1031 net2469 net2285 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[33\] net658 net2622
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[33\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[73\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[73\]
+ net2842 i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_a21oi_1_A1_Y net2834 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q net3268 VGND VPWR i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[254\] clknet_leaf_92_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[421\]_sg13g2_o21ai_1_A1 net3091 VPWR i_snitch.i_snitch_regfile.mem\[421\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[421\] net2810 sg13g2_o21ai_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2610 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ net2919 sg13g2_a221oi_1
XFILLER_103_708 VPWR VGND sg13g2_decap_8
XFILLER_89_909 VPWR VGND sg13g2_decap_8
XFILLER_6_692 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_5_clk clknet_5_0__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A
+ VPWR VGND i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N
+ sg13g2_nand2b_2
XFILLER_38_0 VPWR VGND sg13g2_fill_2
XFILLER_97_964 VPWR VGND sg13g2_decap_8
Xfanout2890 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1_X
+ net2890 VPWR VGND sg13g2_buf_8
XFILLER_84_647 VPWR VGND sg13g2_fill_1
XFILLER_49_390 VPWR VGND sg13g2_fill_2
XFILLER_52_500 VPWR VGND sg13g2_decap_8
XFILLER_37_563 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_fill_1
XFILLER_80_875 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]
+ net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_21_920 VPWR VGND sg13g2_decap_4
XFILLER_33_27 VPWR VGND sg13g2_fill_2
XFILLER_33_49 VPWR VGND sg13g2_fill_2
XFILLER_33_791 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[0\]_sg13g2_nor2_1_A net527 net2732 shift_reg_q\[0\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[2\]_sg13g2_nor2_1_B i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_A i_snitch.pc_d\[2\]
+ i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_Y VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_nor2_1_B
+ net2961 net2954 i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_B1 VPWR VGND
+ sg13g2_nor2_1
XFILLER_106_502 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]_sg13g2_dfrbpq_1_Q
+ net3199 VGND VPWR net604 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net1037 net2452 net2247 VPWR VGND sg13g2_a22oi_1
XFILLER_106_579 VPWR VGND sg13g2_decap_8
XFILLER_88_931 VPWR VGND sg13g2_decap_8
XFILLER_0_835 VPWR VGND sg13g2_decap_8
XFILLER_102_752 VPWR VGND sg13g2_fill_2
XFILLER_102_741 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C
+ VPWR VGND sg13g2_a21o_1
XFILLER_101_273 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2394 net1000 net2469 net2253 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_56_883 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q net3287 VGND VPWR i_snitch.i_snitch_regfile.mem\[274\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[274\] clknet_leaf_93_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[93\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[93\]
+ net2843 i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
XFILLER_15_235 VPWR VGND sg13g2_fill_2
XFILLER_16_758 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2549 VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ VGND net2715 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ sg13g2_o21ai_1
XFILLER_7_467 VPWR VGND sg13g2_decap_8
XFILLER_7_445 VPWR VGND sg13g2_decap_4
XFILLER_99_42 VPWR VGND sg13g2_decap_8
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X
+ net3163 i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nor2b_1_B_N_Y VPWR VGND sg13g2_and3_2
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[409\] clknet_leaf_115_clk sg13g2_dfrbpq_1
Xrsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[16\]_sg13g2_dfrbpq_1_Q_D
+ net951 VGND sg13g2_inv_1
Xdata_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y
+ i_snitch.gpr_waddr\[4\] data_pvalid_sg13g2_nor2b_1_B_N_Y VPWR VGND sg13g2_nand2_1
XFILLER_79_986 VPWR VGND sg13g2_decap_8
XFILLER_94_945 VPWR VGND sg13g2_decap_8
XFILLER_93_400 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]
+ net3165 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2699 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_1 i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_1_Y
+ net2994 i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_nand2b_1_A_N_Y net3022 i_snitch.i_snitch_regfile.mem\[52\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_53_308 VPWR VGND sg13g2_decap_4
XFILLER_47_872 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_0_1017 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[36\]_sg13g2_nor3_1_A net1379 net2767 i_snitch.sb_d\[1\]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[36\]_sg13g2_nor3_1_A_Y VPWR VGND sg13g2_nor3_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A_Y
+ sg13g2_nand4_1
XFILLER_0_1028 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_q\[10\]_sg13g2_dfrbpq_1_Q net3255 VGND VPWR i_snitch.sb_d\[10\] i_snitch.sb_q\[10\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y net2512
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_21_205 VPWR VGND sg13g2_decap_8
XFILLER_22_728 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2631 VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2636 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xhold902 i_snitch.i_snitch_regfile.mem\[75\] VPWR VGND net934 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2390 net793 net2677 net3041 VPWR VGND sg13g2_a22oi_1
Xhold913 data_pdata\[25\] VPWR VGND net945 sg13g2_dlygate4sd3_1
XFILLER_89_706 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y
+ i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_X i_snitch.pc_d\[15\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D_Y
+ VPWR VGND sg13g2_nor4_1
Xhold935 data_pdata\[15\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net967 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[511\]
+ net2802 i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xhold924 i_snitch.i_snitch_regfile.mem\[497\] VPWR VGND net956 sg13g2_dlygate4sd3_1
XFILLER_7_990 VPWR VGND sg13g2_decap_8
Xhold946 i_snitch.i_snitch_regfile.mem\[51\] VPWR VGND net978 sg13g2_dlygate4sd3_1
Xhold968 i_snitch.i_snitch_regfile.mem\[379\] VPWR VGND net1000 sg13g2_dlygate4sd3_1
Xhold957 i_snitch.i_snitch_regfile.mem\[274\] VPWR VGND net989 sg13g2_dlygate4sd3_1
Xhold979 i_snitch.i_snitch_regfile.mem\[60\] VPWR VGND net1011 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2595 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A
+ sg13g2_a21oi_1
XFILLER_88_249 VPWR VGND sg13g2_decap_4
XFILLER_88_227 VPWR VGND sg13g2_fill_2
XFILLER_9_1020 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q net3277 VGND VPWR i_snitch.i_snitch_regfile.mem\[294\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[294\] clknet_leaf_76_clk sg13g2_dfrbpq_1
XFILLER_97_772 VPWR VGND sg13g2_fill_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_97_783 VPWR VGND sg13g2_fill_2
XFILLER_85_934 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] net3178 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_56_146 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net3039
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
XFILLER_56_157 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2735 shift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2
+ shift_reg_q\[24\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[24\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_53_842 VPWR VGND sg13g2_decap_8
XFILLER_25_511 VPWR VGND sg13g2_decap_8
XFILLER_53_864 VPWR VGND sg13g2_fill_1
XFILLER_25_555 VPWR VGND sg13g2_decap_8
XFILLER_100_21 VPWR VGND sg13g2_decap_8
XFILLER_80_683 VPWR VGND sg13g2_decap_8
XFILLER_52_396 VPWR VGND sg13g2_fill_1
XFILLER_52_385 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[466\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_40_525 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A_Y net2840 i_snitch.i_snitch_regfile.mem\[327\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[359\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_100_98 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q net3288 VGND VPWR i_snitch.i_snitch_regfile.mem\[429\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[429\] clknet_leaf_87_clk sg13g2_dfrbpq_1
XFILLER_60_69 VPWR VGND sg13g2_fill_1
XFILLER_5_949 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[218\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[218\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net1092 net2439 net2254 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]
+ net3166 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_106_343 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[113\] clknet_leaf_82_clk sg13g2_dfrbpq_1
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X
+ i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2 net2507 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y
+ VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X
+ sg13g2_nand2b_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2422 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_0_632 VPWR VGND sg13g2_decap_8
XFILLER_102_571 VPWR VGND sg13g2_decap_4
XFILLER_94_219 VPWR VGND sg13g2_fill_1
XFILLER_75_400 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_nand3_1
XFILLER_36_809 VPWR VGND sg13g2_fill_1
XFILLER_91_926 VPWR VGND sg13g2_decap_8
XFILLER_78_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_179 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[12\]_sg13g2_dfrbpq_1_Q net3230 VGND VPWR net549 shift_reg_q\[12\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_71_650 VPWR VGND sg13g2_fill_2
Xi_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_B1 VPWR i_snitch.sb_d\[3\]
+ VGND i_snitch.sb_d\[3\]_sg13g2_o21ai_1_Y_A1 net2293 sg13g2_o21ai_1
XFILLER_43_341 VPWR VGND sg13g2_decap_4
XFILLER_44_897 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[109\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[109\]
+ net2804 sg13g2_o21ai_1
XFILLER_31_503 VPWR VGND sg13g2_decap_8
Xuio_out_sg13g2_buf_1_X_1 i_req_register.data_o\[43\] net14 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_102_1028 VPWR VGND sg13g2_fill_1
XFILLER_102_1017 VPWR VGND sg13g2_decap_8
XFILLER_79_7 VPWR VGND sg13g2_fill_2
XFILLER_7_220 VPWR VGND sg13g2_fill_2
XFILLER_11_271 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[481\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[481\]
+ net2950 sg13g2_o21ai_1
XFILLER_8_776 VPWR VGND sg13g2_fill_2
XFILLER_7_286 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B_sg13g2_o21ai_1_Y
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B
+ sg13g2_o21ai_1
XFILLER_3_492 VPWR VGND sg13g2_decap_8
XFILLER_79_783 VPWR VGND sg13g2_fill_1
XFILLER_66_411 VPWR VGND sg13g2_fill_2
XFILLER_94_753 VPWR VGND sg13g2_fill_2
XFILLER_15_2 VPWR VGND sg13g2_fill_1
XFILLER_38_135 VPWR VGND sg13g2_decap_4
XFILLER_93_252 VPWR VGND sg13g2_fill_1
XFILLER_82_937 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_fill_1
XFILLER_38_168 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1
+ net89 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[449\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[449\] clknet_leaf_75_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[238\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[238\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net835 net2688 net2876 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]
+ net3173 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_35_886 VPWR VGND sg13g2_decap_8
XFILLER_35_897 VPWR VGND sg13g2_fill_2
XFILLER_14_29 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1
+ net2722 i_snitch.inst_addr_o\[11\] i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q net3217 VGND VPWR i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[133\] clknet_leaf_3_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_B
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1
+ net2600 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_30_28 VPWR VGND sg13g2_fill_2
Xhold710 i_snitch.i_snitch_regfile.mem\[448\] VPWR VGND net742 sg13g2_dlygate4sd3_1
Xhold721 i_snitch.i_snitch_regfile.mem\[374\] VPWR VGND net753 sg13g2_dlygate4sd3_1
Xhold743 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\] VPWR
+ VGND net775 sg13g2_dlygate4sd3_1
Xhold732 i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_Y VPWR VGND net764 sg13g2_dlygate4sd3_1
XFILLER_2_908 VPWR VGND sg13g2_decap_8
Xhold754 i_snitch.i_snitch_regfile.mem\[326\] VPWR VGND net786 sg13g2_dlygate4sd3_1
XFILLER_104_858 VPWR VGND sg13g2_decap_8
Xhold776 i_snitch.i_snitch_regfile.mem\[216\] VPWR VGND net808 sg13g2_dlygate4sd3_1
Xhold765 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\] VPWR
+ VGND net797 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[333\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[333\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[333\] net2951 VPWR VGND sg13g2_nand2_1
Xhold787 data_pdata\[26\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net819 sg13g2_dlygate4sd3_1
XFILLER_103_357 VPWR VGND sg13g2_decap_8
Xhold798 i_snitch.i_snitch_regfile.mem\[57\] VPWR VGND net830 sg13g2_dlygate4sd3_1
XFILLER_39_37 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_2
Xi_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0 net3137 i_snitch.i_snitch_regfile.mem\[404\]
+ i_snitch.i_snitch_regfile.mem\[436\] i_snitch.i_snitch_regfile.mem\[468\] i_snitch.i_snitch_regfile.mem\[500\]
+ net3111 i_snitch.i_snitch_regfile.mem\[404\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xshift_reg_q\[0\]_sg13g2_a22oi_1_A1 uio_out_sg13g2_inv_1_Y_3_A shift_reg_q\[0\]_sg13g2_a22oi_1_A1_B1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_1_X
+ cnt_q\[2\]_sg13g2_a22oi_1_B2_A2 shift_reg_q\[0\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y net2723
+ i_snitch.inst_addr_o\[19\] VPWR VGND sg13g2_a22oi_1
XFILLER_69_282 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y
+ i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a21oi_1_A1_A2 i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_mux4_1_A0_1_X
+ VPWR VGND sg13g2_nand2b_1
XFILLER_73_926 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.gpr_waddr\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y
+ i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_2
XFILLER_26_831 VPWR VGND sg13g2_fill_1
XFILLER_81_970 VPWR VGND sg13g2_decap_8
Xdata_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y
+ net2683 data_pdata\[20\]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y VPWR VGND sg13g2_nand2_2
XFILLER_44_149 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[284\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_13_525 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q
+ net3185 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[338\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[338\] VGND sg13g2_inv_1
XFILLER_40_333 VPWR VGND sg13g2_fill_1
XFILLER_41_889 VPWR VGND sg13g2_fill_1
XFILLER_40_388 VPWR VGND sg13g2_decap_8
XFILLER_4_212 VPWR VGND sg13g2_decap_8
XFILLER_106_140 VPWR VGND sg13g2_decap_8
XFILLER_105_0 VPWR VGND sg13g2_decap_8
Xdata_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1 net2683 VPWR data_pdata\[30\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[30\]_sg13g2_a21oi_1_A2_Y net3069 sg13g2_o21ai_1
XFILLER_1_930 VPWR VGND sg13g2_decap_8
XFILLER_20_72 VPWR VGND sg13g2_fill_2
XFILLER_96_21 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y
+ net3087 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q net3262 VGND VPWR i_snitch.i_snitch_regfile.mem\[469\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[469\] clknet_leaf_114_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[430\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[430\]
+ net3018 i_snitch.i_snitch_regfile.mem\[430\]_sg13g2_a21oi_1_A1_Y net2988 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[452\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[452\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[452\] net2947 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ net2599 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[488\]_sg13g2_dfrbpq_1_Q_D VGND net2279 net2365
+ sg13g2_o21ai_1
XFILLER_75_274 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q net3213 VGND VPWR i_snitch.i_snitch_regfile.mem\[153\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[153\] clknet_leaf_116_clk sg13g2_dfrbpq_1
XFILLER_90_244 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A_Y net2947 i_snitch.i_snitch_regfile.mem\[71\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2940 sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[43\]_sg13g2_inv_1_A
+ net844 i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_A2 VPWR VGND sg13g2_inv_4
XFILLER_32_856 VPWR VGND sg13g2_decap_8
XFILLER_32_889 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2379
+ sg13g2_o21ai_1
XFILLER_8_540 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor3_1
XFILLER_6_63 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_99_867 VPWR VGND sg13g2_decap_8
XFILLER_98_366 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[59\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_6_1012 VPWR VGND sg13g2_decap_8
XFILLER_100_338 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2
+ net2716 i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_79_591 VPWR VGND sg13g2_fill_2
Xdata_pdata\[29\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2682 VPWR data_pdata\[29\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[29\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
XFILLER_39_444 VPWR VGND sg13g2_decap_4
XFILLER_66_252 VPWR VGND sg13g2_fill_2
Xrebuffer35 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A
+ net67 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1
+ net2752 net3086 i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[262\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xrebuffer46 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B
+ net78 VPWR VGND sg13g2_buf_1
Xrebuffer24 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1 net56 VPWR VGND sg13g2_buf_1
Xrebuffer13 i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ net45 VPWR VGND sg13g2_buf_8
XFILLER_66_285 VPWR VGND sg13g2_fill_1
XFILLER_27_628 VPWR VGND sg13g2_fill_1
Xrebuffer57 net2609 net89 VPWR VGND sg13g2_buf_1
Xrebuffer68 net2537 net100 VPWR VGND sg13g2_buf_1
Xrebuffer79 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ net111 VPWR VGND sg13g2_buf_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]_sg13g2_nor2_1_B
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[15\]
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.inst_addr_o\[28\]
+ net2523 VPWR VGND sg13g2_xnor2_1
XFILLER_54_447 VPWR VGND sg13g2_fill_2
XFILLER_19_190 VPWR VGND sg13g2_fill_1
XFILLER_81_288 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[468\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[468\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_dfrbpq_1_Q_D VGND net2265 net2357
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2407 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2468 net674 i_snitch.i_snitch_regfile.mem\[389\]_sg13g2_dfrbpq_1_Q_D net2387
+ sg13g2_a221oi_1
Xi_snitch.consec_pc\[0\]_sg13g2_a22oi_1_A1 i_snitch.consec_pc\[0\]_sg13g2_a22oi_1_A1_Y
+ net2628 net49 net2755 i_snitch.consec_pc\[0\] VPWR VGND sg13g2_a22oi_1
XFILLER_50_631 VPWR VGND sg13g2_decap_8
XFILLER_34_182 VPWR VGND sg13g2_decap_4
XFILLER_35_694 VPWR VGND sg13g2_decap_4
XFILLER_10_506 VPWR VGND sg13g2_decap_4
XFILLER_23_889 VPWR VGND sg13g2_decap_8
XFILLER_50_697 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q net3275 VGND VPWR i_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[489\] clknet_leaf_105_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[278\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2325 net944 net2652 net2893 VPWR VGND sg13g2_a22oi_1
XFILLER_2_705 VPWR VGND sg13g2_decap_8
Xfanout2708 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X
+ net2708 VPWR VGND sg13g2_buf_8
Xhold562 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\] VPWR
+ VGND net594 sg13g2_dlygate4sd3_1
Xhold551 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net583 sg13g2_dlygate4sd3_1
XFILLER_9_7 VPWR VGND sg13g2_decap_8
Xhold540 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net572 sg13g2_dlygate4sd3_1
Xhold573 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[1\] VPWR
+ VGND net605 sg13g2_dlygate4sd3_1
XFILLER_89_355 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xfanout2719 net2721 net2719 VPWR VGND sg13g2_buf_8
Xhold584 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\] VPWR
+ VGND net616 sg13g2_dlygate4sd3_1
Xhold595 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\] VPWR
+ VGND net627 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q net3296 VGND VPWR i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[173\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_106_42 VPWR VGND sg13g2_decap_8
XFILLER_103_154 VPWR VGND sg13g2_decap_8
XFILLER_100_861 VPWR VGND sg13g2_decap_8
XFILLER_85_550 VPWR VGND sg13g2_decap_4
Xhold1240 rsp_data_q\[23\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1272
+ sg13g2_dlygate4sd3_1
XFILLER_57_263 VPWR VGND sg13g2_decap_8
Xhold1251 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] VPWR
+ VGND net1283 sg13g2_dlygate4sd3_1
Xhold1262 rsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1294
+ sg13g2_dlygate4sd3_1
XFILLER_72_200 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0 net3123 i_snitch.i_snitch_regfile.mem\[287\]
+ i_snitch.i_snitch_regfile.mem\[319\] i_snitch.i_snitch_regfile.mem\[351\] i_snitch.i_snitch_regfile.mem\[383\]
+ net3113 i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xhold1284 i_snitch.i_snitch_regfile.mem\[289\] VPWR VGND net1316 sg13g2_dlygate4sd3_1
Xhold1273 i_snitch.i_snitch_regfile.mem\[100\] VPWR VGND net1305 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y
+ VPWR VGND sg13g2_nor3_2
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A_sg13g2_or2_1_X
+ VGND VPWR data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A
+ net3141 net3144 sg13g2_or2_1
Xhold1295 i_snitch.i_snitch_regfile.mem\[227\] VPWR VGND net1327 sg13g2_dlygate4sd3_1
XFILLER_54_992 VPWR VGND sg13g2_fill_2
XFILLER_72_299 VPWR VGND sg13g2_fill_2
Xheichips25_snitch_wrapper_28 VPWR VGND uio_oe[4] sg13g2_tiehi
XFILLER_13_377 VPWR VGND sg13g2_decap_8
XFILLER_14_889 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q net3316 VGND VPWR i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[308\] clknet_leaf_66_clk sg13g2_dfrbpq_1
XFILLER_9_326 VPWR VGND sg13g2_fill_1
XFILLER_99_119 VPWR VGND sg13g2_decap_8
XFILLER_96_859 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[502\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2365
+ sg13g2_o21ai_1
XFILLER_49_731 VPWR VGND sg13g2_fill_2
XFILLER_95_369 VPWR VGND sg13g2_fill_2
XFILLER_76_561 VPWR VGND sg13g2_fill_1
XFILLER_49_786 VPWR VGND sg13g2_decap_8
XFILLER_0_292 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
XFILLER_37_926 VPWR VGND sg13g2_fill_2
XFILLER_48_285 VPWR VGND sg13g2_fill_1
XFILLER_36_425 VPWR VGND sg13g2_fill_1
XFILLER_63_244 VPWR VGND sg13g2_decap_4
XFILLER_36_469 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2 VGND
+ VPWR net2965 i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1_X i_snitch.i_snitch_regfile.mem\[396\]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[332\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_45_970 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[298\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[298\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2431 net2283 net2317 net1257 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2478 i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2457 net2856 i_snitch.i_snitch_regfile.mem\[483\]_sg13g2_dfrbpq_1_Q_D net2910
+ sg13g2_a221oi_1
XFILLER_17_694 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ net2415 sg13g2_a21oi_1
Xdata_pdata\[3\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C net3149 data_pdata\[11\]_sg13g2_nor2b_1_A_Y
+ data_pdata\[3\]_sg13g2_nor2_1_B_Y data_pdata\[3\]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_60_973 VPWR VGND sg13g2_fill_1
XFILLER_20_804 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[104\]_sg13g2_o21ai_1_A1_Y net3090 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[392\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[360\]_sg13g2_o21ai_1_A1 net2971 VPWR i_snitch.i_snitch_regfile.mem\[360\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[360\] net2808 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q net3279 VGND VPWR i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[193\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_68_0 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ net2498 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X VPWR
+ VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[299\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[299\]
+ net3021 i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_a21oi_1_A1_Y net2990 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[324\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[324\] VGND sg13g2_inv_1
XFILLER_87_804 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[41\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[41\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_59_517 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[472\]_sg13g2_dfrbpq_1_Q_D VGND net2256 net2378
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[459\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_nand2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[459\] net2953 VPWR VGND sg13g2_nand2_1
XFILLER_28_904 VPWR VGND sg13g2_fill_2
XFILLER_39_252 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[328\]_sg13g2_dfrbpq_1_Q net3307 VGND VPWR i_snitch.i_snitch_regfile.mem\[328\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[328\] clknet_leaf_74_clk sg13g2_dfrbpq_1
XFILLER_27_403 VPWR VGND sg13g2_decap_8
XFILLER_27_458 VPWR VGND sg13g2_fill_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ net2720 VPWR VGND sg13g2_nand2_1
XFILLER_70_737 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1 VGND i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_55_789 VPWR VGND sg13g2_fill_2
XFILLER_54_288 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[117\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2449 net2269 net2409 net1204 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[142\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2274
+ net2446 VPWR VGND sg13g2_nand2_1
XFILLER_22_185 VPWR VGND sg13g2_decap_8
XFILLER_7_808 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[16\]_sg13g2_a22oi_1_A1 shift_reg_q\[16\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_mux2_1_A1_1_X
+ net3057 net3047 net546 VPWR VGND sg13g2_a22oi_1
XFILLER_105_931 VPWR VGND sg13g2_decap_8
Xfanout3228 net3229 net3228 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[374\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[278\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[342\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2847
+ sg13g2_a221oi_1
Xfanout3206 net3208 net3206 VPWR VGND sg13g2_buf_8
Xfanout3217 net3225 net3217 VPWR VGND sg13g2_buf_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
Xfanout3239 net3249 net3239 VPWR VGND sg13g2_buf_8
Xfanout2527 net2528 net2527 VPWR VGND sg13g2_buf_8
Xfanout2516 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y
+ net2516 VPWR VGND sg13g2_buf_1
XFILLER_7_4 VPWR VGND sg13g2_decap_8
Xfanout2505 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y
+ net2505 VPWR VGND sg13g2_buf_8
Xfanout2538 net2539 net2538 VPWR VGND sg13g2_buf_8
Xfanout2549 net2550 net2549 VPWR VGND sg13g2_buf_8
XFILLER_81_1026 VPWR VGND sg13g2_fill_2
Xhold392 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\] VPWR
+ VGND net424 sg13g2_dlygate4sd3_1
XFILLER_104_496 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D
+ VPWR VGND sg13g2_nor3_1
XFILLER_93_807 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A
+ i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B i_snitch.i_snitch_lsu.handshake_pending_d
+ VPWR VGND sg13g2_nor2_1
XFILLER_58_561 VPWR VGND sg13g2_decap_8
XFILLER_86_881 VPWR VGND sg13g2_decap_8
XFILLER_73_520 VPWR VGND sg13g2_fill_1
XFILLER_58_572 VPWR VGND sg13g2_fill_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B net2795
+ i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_46_767 VPWR VGND sg13g2_decap_4
XFILLER_18_447 VPWR VGND sg13g2_fill_2
Xhold1070 i_snitch.i_snitch_regfile.mem\[358\] VPWR VGND net1102 sg13g2_dlygate4sd3_1
Xhold1092 i_snitch.i_snitch_regfile.mem\[46\] VPWR VGND net1124 sg13g2_dlygate4sd3_1
Xhold1081 i_snitch.i_snitch_regfile.mem\[198\] VPWR VGND net1113 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_dfrbpq_1_Q_D VGND net2243 net2363
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net950 net2494 net1303 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2724 i_snitch.inst_addr_o\[12\] sg13g2_a21oi_2
XFILLER_14_664 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ sg13g2_nand2b_2
Xi_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[403\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net3038
+ net2673 VPWR VGND sg13g2_nand2_1
XFILLER_41_461 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q net3270 VGND VPWR i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[61\] clknet_leaf_94_clk sg13g2_dfrbpq_1
Xreq_data_valid_sg13g2_o21ai_1_Y req_data_valid_sg13g2_o21ai_1_Y_B1 VPWR req_data_valid
+ VGND net3053 i_req_register.data_o\[5\]_sg13g2_inv_1_A_Y sg13g2_o21ai_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y
+ VGND net3148 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X
+ sg13g2_o21ai_1
Xrebuffer4 net35 net36 VPWR VGND sg13g2_buf_1
Xi_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A VPWR
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y VGND sg13g2_inv_1
XFILLER_5_340 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[454\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[454\] VGND sg13g2_inv_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2600 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_6_885 VPWR VGND sg13g2_fill_2
XFILLER_6_874 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q net3263 VGND VPWR i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[348\] clknet_leaf_97_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[507\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2854
+ net2658 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[173\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2444 VPWR VGND sg13g2_nand2_1
XFILLER_96_656 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2352 net738 net2686 net2887 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_B1 VPWR
+ i_snitch.sb_d\[10\] VGND net2292 i_snitch.sb_d\[10\]_sg13g2_o21ai_1_Y_A2 sg13g2_o21ai_1
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_56_509 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[320\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2400
+ sg13g2_o21ai_1
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[57\]_sg13g2_o21ai_1_A1 net3004 VPWR i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[57\] net2977 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1 net3120 i_snitch.i_snitch_regfile.mem\[131\]
+ i_snitch.i_snitch_regfile.mem\[163\] i_snitch.i_snitch_regfile.mem\[195\] i_snitch.i_snitch_regfile.mem\[227\]
+ net3101 i_snitch.i_snitch_regfile.mem\[131\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net43 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_36_233 VPWR VGND sg13g2_decap_4
XFILLER_37_778 VPWR VGND sg13g2_fill_2
XFILLER_52_748 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[277\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2670 VPWR VGND sg13g2_nand2_1
XFILLER_20_634 VPWR VGND sg13g2_fill_1
XFILLER_32_483 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ VGND net2750 net2589 sg13g2_o21ai_1
XFILLER_20_678 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2798
+ net2693 VPWR VGND sg13g2_nand2_1
XFILLER_106_706 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2
+ net3009 sg13g2_a21oi_2
Xdata_pdata\[2\]_sg13g2_dfrbpq_1_Q net3202 VGND VPWR net687 data_pdata\[2\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_105_238 VPWR VGND sg13g2_decap_8
XFILLER_102_912 VPWR VGND sg13g2_decap_8
XFILLER_59_303 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2510 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2 net2831
+ VPWR i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.i_snitch_regfile.mem\[117\]_sg13g2_nor2_1_A_1_Y i_snitch.i_snitch_regfile.mem\[53\]_sg13g2_a22oi_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_102_989 VPWR VGND sg13g2_decap_8
XFILLER_47_509 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[434\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2864
+ net2675 VPWR VGND sg13g2_nand2_1
XFILLER_74_339 VPWR VGND sg13g2_decap_8
XFILLER_68_870 VPWR VGND sg13g2_fill_2
XFILLER_103_21 VPWR VGND sg13g2_decap_8
XFILLER_83_851 VPWR VGND sg13g2_decap_8
XFILLER_82_350 VPWR VGND sg13g2_fill_2
XFILLER_43_715 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[81\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[81\] clknet_leaf_82_clk sg13g2_dfrbpq_1
XFILLER_42_203 VPWR VGND sg13g2_fill_2
XFILLER_103_98 VPWR VGND sg13g2_decap_8
XFILLER_27_299 VPWR VGND sg13g2_decap_8
XFILLER_51_792 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q net3286 VGND VPWR i_snitch.i_snitch_regfile.mem\[368\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[368\] clknet_leaf_86_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y
+ VGND VPWR net2550 i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
XFILLER_6_126 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[12\] net1049 net2917 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[157\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[157\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2351 net1098 net2446 net2250 VPWR VGND sg13g2_a22oi_1
XFILLER_3_822 VPWR VGND sg13g2_decap_8
Xfanout3003 net3011 net3003 VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2552 VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1
+ VGND net2715 i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ sg13g2_o21ai_1
Xfanout3036 net3037 net3036 VPWR VGND sg13g2_buf_1
Xfanout2302 net2311 net2302 VPWR VGND sg13g2_buf_8
Xfanout3025 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y
+ net3025 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1 net3001 i_snitch.i_snitch_regfile.mem\[133\]
+ i_snitch.i_snitch_regfile.mem\[165\] i_snitch.i_snitch_regfile.mem\[197\] i_snitch.i_snitch_regfile.mem\[229\]
+ net2974 i_snitch.i_snitch_regfile.mem\[133\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xfanout3014 net3015 net3014 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[77\]_sg13g2_o21ai_1_A1 net2988 VPWR i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[77\] net3017 sg13g2_o21ai_1
Xfanout3058 net3059 net3058 VPWR VGND sg13g2_buf_8
Xfanout2313 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ net2313 VPWR VGND sg13g2_buf_1
Xfanout3047 cnt_q\[2\]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X net3047 VPWR VGND sg13g2_buf_2
Xfanout2335 i_snitch.sb_d\[6\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2335 VPWR VGND sg13g2_buf_8
Xfanout2324 net2327 net2324 VPWR VGND sg13g2_buf_8
Xfanout3069 i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_nand2b_1_B_Y net3069 VPWR
+ VGND sg13g2_buf_8
Xfanout2357 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ net2357 VPWR VGND sg13g2_buf_8
Xfanout2368 net2370 net2368 VPWR VGND sg13g2_buf_8
XFILLER_3_899 VPWR VGND sg13g2_decap_8
Xfanout2346 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y
+ net2346 VPWR VGND sg13g2_buf_8
Xfanout2379 net2380 net2379 VPWR VGND sg13g2_buf_8
XFILLER_38_509 VPWR VGND sg13g2_decap_4
XFILLER_78_689 VPWR VGND sg13g2_decap_8
Xshift_reg_q\[14\]_sg13g2_nor2_1_A net486 net2733 shift_reg_q\[14\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_19_712 VPWR VGND sg13g2_decap_4
XFILLER_19_734 VPWR VGND sg13g2_fill_1
XFILLER_74_862 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2700 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_33_214 VPWR VGND sg13g2_decap_4
Xdata_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1 data_pdata\[11\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y
+ data_pdata\[27\]_sg13g2_nand2b_1_B_Y net3151 data_pdata\[19\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[11\]_sg13g2_nand2b_1_B_Y VPWR VGND sg13g2_a22oi_1
XFILLER_21_409 VPWR VGND sg13g2_fill_1
XFILLER_33_269 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[108\]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.inst_addr_o\[28\]_sg13g2_dfrbpq_1_Q net3305 VGND VPWR i_snitch.pc_d\[28\]
+ i_snitch.inst_addr_o\[28\] clknet_leaf_51_clk sg13g2_dfrbpq_2
XFILLER_105_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2470
+ net2513 net2901 net2881 VPWR VGND sg13g2_a22oi_1
XFILLER_97_943 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X
+ net3072 i_snitch.sb_q\[12\] i_snitch.sb_q\[13\] i_snitch.sb_q\[14\] i_snitch.sb_q\[15\]
+ net3071 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_mux4_1
XFILLER_69_678 VPWR VGND sg13g2_decap_4
XFILLER_68_144 VPWR VGND sg13g2_fill_2
Xfanout2891 net2896 net2891 VPWR VGND sg13g2_buf_8
Xfanout2880 net2884 net2880 VPWR VGND sg13g2_buf_8
XFILLER_96_475 VPWR VGND sg13g2_fill_1
XFILLER_84_637 VPWR VGND sg13g2_decap_4
XFILLER_92_670 VPWR VGND sg13g2_decap_8
XFILLER_83_158 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2458
+ net2244 net2649 net2858 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q net3219 VGND VPWR i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[388\] clknet_leaf_14_clk sg13g2_dfrbpq_1
Xi_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[4\]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[177\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[177\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2345 net727 net2664 net2775 VPWR VGND sg13g2_a22oi_1
Xi_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 net2627 net2757 i_snitch.pc_d\[25\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1 net2999 i_snitch.i_snitch_regfile.mem\[135\]
+ i_snitch.i_snitch_regfile.mem\[167\] i_snitch.i_snitch_regfile.mem\[199\] i_snitch.i_snitch_regfile.mem\[231\]
+ net2973 i_snitch.i_snitch_regfile.mem\[135\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_20_420 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1 net2832 VPWR i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[97\] net3026 sg13g2_o21ai_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X
+ i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B
+ VPWR VGND sg13g2_xor2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2706 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1
+ net2614 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_nor2_1_Y
+ net2568 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_4_619 VPWR VGND sg13g2_fill_1
XFILLER_106_558 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2934 i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[55\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
XFILLER_88_910 VPWR VGND sg13g2_decap_8
XFILLER_0_814 VPWR VGND sg13g2_decap_8
XFILLER_102_720 VPWR VGND sg13g2_fill_2
XFILLER_99_280 VPWR VGND sg13g2_decap_8
XFILLER_87_420 VPWR VGND sg13g2_fill_2
XFILLER_88_987 VPWR VGND sg13g2_decap_8
XFILLER_87_442 VPWR VGND sg13g2_decap_4
Xshift_reg_q\[27\]_sg13g2_nor2_1_A net614 net2737 shift_reg_q\[27\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_102_786 VPWR VGND sg13g2_decap_8
XFILLER_101_252 VPWR VGND sg13g2_decap_8
XFILLER_87_486 VPWR VGND sg13g2_fill_1
XFILLER_87_475 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q net3298 VGND VPWR i_snitch.i_snitch_regfile.mem\[207\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[207\] clknet_leaf_81_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[496\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2858
+ net2667 VPWR VGND sg13g2_nand2_1
XFILLER_56_862 VPWR VGND sg13g2_fill_2
XFILLER_28_553 VPWR VGND sg13g2_fill_2
XFILLER_83_692 VPWR VGND sg13g2_decap_8
XFILLER_71_843 VPWR VGND sg13g2_decap_4
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_12_965 VPWR VGND sg13g2_fill_1
XFILLER_7_413 VPWR VGND sg13g2_fill_1
XFILLER_99_21 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_inv_1_Y
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X
+ VGND sg13g2_inv_1
XFILLER_8_969 VPWR VGND sg13g2_decap_8
XFILLER_87_1021 VPWR VGND sg13g2_decap_8
XFILLER_99_98 VPWR VGND sg13g2_decap_8
XFILLER_3_630 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2713 i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B_X
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2786
+ net2650 VPWR VGND sg13g2_nand2_1
XFILLER_3_685 VPWR VGND sg13g2_fill_2
XFILLER_3_674 VPWR VGND sg13g2_decap_8
XFILLER_79_965 VPWR VGND sg13g2_decap_8
XFILLER_94_924 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[503\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2370 net784 net2647 net2857 VPWR VGND sg13g2_a22oi_1
XFILLER_38_306 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B
+ VGND net2594 i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_93_434 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1 net3009 i_snitch.i_snitch_regfile.mem\[137\]
+ i_snitch.i_snitch_regfile.mem\[169\] i_snitch.i_snitch_regfile.mem\[201\] i_snitch.i_snitch_regfile.mem\[233\]
+ net2983 i_snitch.i_snitch_regfile.mem\[137\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_19_531 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ net2577 VPWR VGND sg13g2_a22oi_1
XFILLER_74_670 VPWR VGND sg13g2_fill_2
XFILLER_62_810 VPWR VGND sg13g2_fill_2
XFILLER_47_884 VPWR VGND sg13g2_fill_1
XFILLER_47_862 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_fill_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_80_139 VPWR VGND sg13g2_decap_4
XFILLER_74_681 VPWR VGND sg13g2_decap_4
XFILLER_0_98 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1046 net2690 net2768 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[45\]_sg13g2_a22oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[77\]_sg13g2_mux2_1_A0_X net3108 net2830 i_snitch.i_snitch_regfile.mem\[45\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_14_280 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[329\] VGND sg13g2_inv_1
XFILLER_30_784 VPWR VGND sg13g2_fill_1
Xstrb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A
+ strb_reg_q\[6\]_sg13g2_nor2_1_A_Y strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D VPWR VGND
+ sg13g2_nor2_1
Xhold903 i_snitch.i_snitch_regfile.mem\[478\] VPWR VGND net935 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.inst_addr_o\[21\]
+ net2526 VPWR VGND sg13g2_xnor2_1
XFILLER_50_0 VPWR VGND sg13g2_fill_1
Xhold925 i_snitch.i_snitch_regfile.mem\[352\] VPWR VGND net957 sg13g2_dlygate4sd3_1
Xhold936 i_snitch.i_snitch_regfile.mem\[210\] VPWR VGND net968 sg13g2_dlygate4sd3_1
Xhold914 data_pdata\[25\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net946 sg13g2_dlygate4sd3_1
XFILLER_89_729 VPWR VGND sg13g2_fill_1
Xhold958 i_snitch.inst_addr_o\[10\] VPWR VGND net990 sg13g2_dlygate4sd3_1
Xhold969 i_snitch.i_snitch_regfile.mem\[495\] VPWR VGND net1001 sg13g2_dlygate4sd3_1
Xhold947 i_snitch.i_snitch_regfile.mem\[241\] VPWR VGND net979 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q net3221 VGND VPWR i_snitch.i_snitch_regfile.mem\[227\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[227\] clknet_leaf_108_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_mux2_1_A1
+ net758 net581 net2240 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[26\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B_sg13g2_and2_1_X net3072
+ net2536 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B VPWR VGND sg13g2_and2_1
Xi_snitch.sb_q\[4\]_sg13g2_dfrbpq_1_Q net3250 VGND VPWR i_snitch.sb_d\[4\] i_snitch.sb_q\[4\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[110\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[46\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_69_453 VPWR VGND sg13g2_decap_4
XFILLER_85_913 VPWR VGND sg13g2_decap_8
XFILLER_69_464 VPWR VGND sg13g2_fill_1
XFILLER_57_604 VPWR VGND sg13g2_fill_1
XFILLER_29_317 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B sg13g2_o21ai_1
XFILLER_72_618 VPWR VGND sg13g2_fill_1
XFILLER_38_873 VPWR VGND sg13g2_fill_1
XFILLER_25_523 VPWR VGND sg13g2_decap_8
XFILLER_38_895 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A
+ VPWR VGND sg13g2_nor3_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C
+ net3076 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[27\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_64_180 VPWR VGND sg13g2_fill_1
XFILLER_52_375 VPWR VGND sg13g2_decap_4
Xdata_pdata\[13\]_sg13g2_nor2b_1_A data_pdata\[13\] net3155 data_pdata\[13\]_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_o21ai_1_A2
+ net2542 VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ VGND net2750 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2
+ sg13g2_o21ai_1
Xdata_pdata\[6\]_sg13g2_mux2_1_A0 data_pdata\[6\] data_pdata\[14\] net3162 data_pdata\[6\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
XFILLER_40_559 VPWR VGND sg13g2_decap_8
Xi_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B net2887 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2
+ net2503 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y VPWR VGND sg13g2_nor3_1
XFILLER_100_77 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y
+ net2637 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y
+ net2719 i_req_arb.data_i\[41\] VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1
+ VPWR VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1
+ net2815 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2698 i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B
+ net2540 sg13g2_a21oi_1
XFILLER_5_928 VPWR VGND sg13g2_decap_8
XFILLER_106_322 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1 net3021 i_snitch.i_snitch_regfile.mem\[139\]
+ i_snitch.i_snitch_regfile.mem\[171\] i_snitch.i_snitch_regfile.mem\[203\] i_snitch.i_snitch_regfile.mem\[235\]
+ net2992 i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_106_399 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2584 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_0_611 VPWR VGND sg13g2_decap_8
XFILLER_88_751 VPWR VGND sg13g2_decap_8
Xstrb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X net2727 net534
+ strb_reg_q\[6\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A VPWR VGND sg13g2_and2_1
XFILLER_0_688 VPWR VGND sg13g2_decap_8
XFILLER_76_946 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[87\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_nand2b_1_A_N_Y
+ net3030 i_snitch.i_snitch_regfile.mem\[87\] VPWR VGND sg13g2_nand2b_1
XFILLER_91_905 VPWR VGND sg13g2_decap_8
XFILLER_29_873 VPWR VGND sg13g2_fill_2
XFILLER_62_106 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_16_501 VPWR VGND sg13g2_decap_8
XFILLER_90_459 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[163\]_sg13g2_nor3_1_A net1309 net2772 i_snitch.sb_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[163\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_71_684 VPWR VGND sg13g2_fill_1
XFILLER_70_150 VPWR VGND sg13g2_decap_4
XFILLER_43_364 VPWR VGND sg13g2_decap_4
XFILLER_16_589 VPWR VGND sg13g2_decap_4
XFILLER_31_559 VPWR VGND sg13g2_fill_2
XFILLER_34_71 VPWR VGND sg13g2_fill_2
XFILLER_34_82 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_C1 net2637 i_snitch.inst_addr_o\[17\]
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ net2724 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q net3328 VGND VPWR i_snitch.i_snitch_regfile.mem\[247\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[247\] clknet_leaf_56_clk sg13g2_dfrbpq_1
Xuio_out_sg13g2_buf_1_X_2 i_req_register.data_o\[44\] net15 VPWR VGND sg13g2_buf_1
Xi_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[14\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y
+ VPWR VGND sg13g2_nand2_2
XFILLER_8_744 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2720 i_snitch.inst_addr_o\[28\] sg13g2_a21oi_2
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B
+ VGND VPWR i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ sg13g2_or2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1
+ net2589 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND sg13g2_a22oi_1
XFILLER_4_983 VPWR VGND sg13g2_decap_8
XFILLER_3_460 VPWR VGND sg13g2_decap_8
XFILLER_61_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A_Y net2828 i_snitch.i_snitch_regfile.mem\[312\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_22_4 VPWR VGND sg13g2_decap_4
XFILLER_67_957 VPWR VGND sg13g2_decap_8
XFILLER_82_916 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.inst_addr_o\[25\] net2523 VPWR VGND sg13g2_nand2_1
XFILLER_66_467 VPWR VGND sg13g2_fill_1
XFILLER_94_798 VPWR VGND sg13g2_fill_1
XFILLER_93_297 VPWR VGND sg13g2_fill_1
XFILLER_81_426 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3061 net1051 net3065 rsp_data_q\[24\] VPWR VGND sg13g2_a22oi_1
XFILLER_47_692 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[345\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_98_0 VPWR VGND sg13g2_decap_8
XFILLER_50_868 VPWR VGND sg13g2_fill_2
XFILLER_50_857 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1
+ net2724 net2965 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_50_879 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C VPWR
+ VGND sg13g2_nor3_2
Xhold700 i_snitch.i_snitch_regfile.mem\[152\] VPWR VGND net732 sg13g2_dlygate4sd3_1
Xhold711 i_snitch.i_snitch_regfile.mem\[342\] VPWR VGND net743 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[85\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[85\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2353 net877 net2452 net2269 VPWR VGND sg13g2_a22oi_1
Xhold744 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net776 sg13g2_dlygate4sd3_1
Xhold733 i_snitch.i_snitch_regfile.mem\[64\] VPWR VGND net765 sg13g2_dlygate4sd3_1
Xhold755 i_snitch.i_snitch_regfile.mem\[267\] VPWR VGND net787 sg13g2_dlygate4sd3_1
Xhold722 data_pdata\[19\] VPWR VGND net754 sg13g2_dlygate4sd3_1
XFILLER_104_837 VPWR VGND sg13g2_decap_8
Xhold777 data_pdata\[16\] VPWR VGND net809 sg13g2_dlygate4sd3_1
Xhold766 data_pdata\[22\] VPWR VGND net798 sg13g2_dlygate4sd3_1
Xhold788 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] VPWR
+ VGND net820 sg13g2_dlygate4sd3_1
XFILLER_103_336 VPWR VGND sg13g2_decap_8
Xhold799 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\] VPWR
+ VGND net831 sg13g2_dlygate4sd3_1
Xi_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1 i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2
+ i_snitch.wake_up_q\[1\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2 net553 VPWR VGND
+ sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[299\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VGND
+ i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_inv_1_A_Y net3020 sg13g2_o21ai_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B
+ sg13g2_or2_1
XFILLER_57_434 VPWR VGND sg13g2_fill_1
XFILLER_55_15 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[267\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q
+ net3246 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_72_437 VPWR VGND sg13g2_fill_2
XFILLER_44_117 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]_sg13g2_dfrbpq_1_Q
+ net3245 VGND VPWR net1050 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[12\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
XFILLER_52_150 VPWR VGND sg13g2_decap_4
XFILLER_13_515 VPWR VGND sg13g2_fill_1
XFILLER_40_301 VPWR VGND sg13g2_fill_1
XFILLER_52_194 VPWR VGND sg13g2_decap_4
XFILLER_40_345 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B_Y
+ net2515 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_4_224 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[254\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_84_1024 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[0\]_sg13g2_dfrbpq_1_Q net3235 VGND
+ VPWR net1332 i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q\[0\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_20_51 VPWR VGND sg13g2_decap_4
XFILLER_4_268 VPWR VGND sg13g2_fill_2
XFILLER_106_196 VPWR VGND sg13g2_decap_8
XFILLER_96_77 VPWR VGND sg13g2_decap_8
XFILLER_49_902 VPWR VGND sg13g2_decap_4
XFILLER_1_986 VPWR VGND sg13g2_decap_8
XFILLER_88_592 VPWR VGND sg13g2_decap_8
XFILLER_76_732 VPWR VGND sg13g2_decap_4
XFILLER_49_946 VPWR VGND sg13g2_fill_2
XFILLER_48_412 VPWR VGND sg13g2_decap_8
XFILLER_64_905 VPWR VGND sg13g2_fill_1
XFILLER_63_404 VPWR VGND sg13g2_decap_8
XFILLER_91_746 VPWR VGND sg13g2_fill_1
XFILLER_63_426 VPWR VGND sg13g2_fill_2
Xrsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ net1184 VGND sg13g2_inv_1
XFILLER_91_768 VPWR VGND sg13g2_decap_8
XFILLER_63_448 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[481\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2
+ net2505 i_snitch.sb_d\[13\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_2
XFILLER_91_1017 VPWR VGND sg13g2_decap_8
XFILLER_90_278 VPWR VGND sg13g2_fill_1
XFILLER_44_673 VPWR VGND sg13g2_fill_2
XFILLER_91_1028 VPWR VGND sg13g2_fill_1
XFILLER_91_7 VPWR VGND sg13g2_decap_8
XFILLER_44_695 VPWR VGND sg13g2_fill_2
XFILLER_43_183 VPWR VGND sg13g2_decap_8
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
XFILLER_40_890 VPWR VGND sg13g2_fill_2
XFILLER_8_585 VPWR VGND sg13g2_fill_2
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_99_846 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q net3302 VGND VPWR i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[287\] clknet_leaf_71_clk sg13g2_dfrbpq_1
XFILLER_100_317 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q
+ net3190 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
XFILLER_94_551 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B
+ VGND i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ sg13g2_o21ai_1
XFILLER_82_702 VPWR VGND sg13g2_fill_2
XFILLER_13_0 VPWR VGND sg13g2_fill_2
XFILLER_94_595 VPWR VGND sg13g2_fill_2
XFILLER_94_584 VPWR VGND sg13g2_fill_2
Xrebuffer14 i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_B
+ net46 VPWR VGND sg13g2_buf_2
Xrebuffer36 net68 net2241 VPWR VGND sg13g2_buf_16
Xrebuffer25 i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1 net57 VPWR VGND sg13g2_buf_1
XFILLER_66_297 VPWR VGND sg13g2_fill_1
XFILLER_66_264 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2408 i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_nor3_1_A_Y net2455 net2765 i_snitch.i_snitch_regfile.mem\[37\]_sg13g2_dfrbpq_1_Q_D
+ net2906 sg13g2_a221oi_1
Xrebuffer69 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ net101 VPWR VGND sg13g2_buf_1
Xrebuffer58 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net90 VPWR VGND sg13g2_buf_1
XFILLER_81_234 VPWR VGND sg13g2_fill_1
XFILLER_70_919 VPWR VGND sg13g2_fill_1
Xrebuffer47 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_X
+ net79 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[97\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[97\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net494 net2409 VPWR VGND sg13g2_nand2_1
Xdata_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[24\]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[24\]_sg13g2_a21oi_1_A2_Y net3068 sg13g2_o21ai_1
XFILLER_62_492 VPWR VGND sg13g2_fill_1
XFILLER_34_172 VPWR VGND sg13g2_fill_1
Xdata_pdata\[26\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1 net2681 VPWR data_pdata\[26\]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y
+ VGND data_pdata\[26\]_sg13g2_nand2b_1_B_Y net3068 sg13g2_o21ai_1
XFILLER_22_367 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[20\]_sg13g2_or2_1_B VGND VPWR i_snitch.pc_d\[20\]_sg13g2_or2_1_B_X
+ i_snitch.pc_d\[20\] i_snitch.inst_addr_o\[20\] sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[102\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[49\]_sg13g2_dfrbpq_1_Q_D VGND net2289 net2363
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[106\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2484 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2468 net3039 i_snitch.i_snitch_regfile.mem\[386\]_sg13g2_dfrbpq_1_Q_D net2911
+ sg13g2_a221oi_1
Xhold530 i_snitch.i_snitch_regfile.mem\[273\] VPWR VGND net562 sg13g2_dlygate4sd3_1
Xfanout2709 net2710 net2709 VPWR VGND sg13g2_buf_8
Xhold563 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net595 sg13g2_dlygate4sd3_1
Xhold552 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\] VPWR
+ VGND net584 sg13g2_dlygate4sd3_1
Xhold541 i_snitch.sb_q\[11\] VPWR VGND net573 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[445\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1 i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[62\]_sg13g2_o21ai_1_A1_Y i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[414\]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y net2954
+ VPWR VGND sg13g2_a22oi_1
XFILLER_103_133 VPWR VGND sg13g2_decap_8
Xhold585 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net617 sg13g2_dlygate4sd3_1
Xhold574 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\] VPWR
+ VGND net606 sg13g2_dlygate4sd3_1
Xhold596 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[40\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net628 sg13g2_dlygate4sd3_1
XFILLER_106_21 VPWR VGND sg13g2_decap_8
XFILLER_89_378 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[367\]_sg13g2_dfrbpq_1_Q_D VGND net2264 net2392
+ sg13g2_o21ai_1
XFILLER_106_98 VPWR VGND sg13g2_decap_8
XFILLER_100_840 VPWR VGND sg13g2_decap_8
XFILLER_85_562 VPWR VGND sg13g2_decap_4
XFILLER_66_58 VPWR VGND sg13g2_decap_8
XFILLER_66_47 VPWR VGND sg13g2_fill_1
Xhold1230 i_snitch.i_snitch_regfile.mem\[410\] VPWR VGND net1262 sg13g2_dlygate4sd3_1
Xhold1241 i_snitch.i_snitch_regfile.mem\[114\] VPWR VGND net1273 sg13g2_dlygate4sd3_1
Xhold1252 i_snitch.i_snitch_regfile.mem\[356\] VPWR VGND net1284 sg13g2_dlygate4sd3_1
Xhold1274 rsp_data_q\[12\] VPWR VGND net1306 sg13g2_dlygate4sd3_1
XFILLER_46_938 VPWR VGND sg13g2_decap_4
XFILLER_45_404 VPWR VGND sg13g2_fill_1
Xhold1285 i_snitch.i_snitch_regfile.mem\[391\] VPWR VGND net1317 sg13g2_dlygate4sd3_1
Xhold1263 i_snitch.i_snitch_regfile.mem\[103\] VPWR VGND net1295 sg13g2_dlygate4sd3_1
XFILLER_18_629 VPWR VGND sg13g2_decap_4
Xhold1296 i_snitch.i_snitch_regfile.mem\[421\] VPWR VGND net1328 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0 net124 i_snitch.i_snitch_regfile.mem\[134\]
+ i_snitch.i_snitch_regfile.mem\[166\] i_snitch.i_snitch_regfile.mem\[198\] i_snitch.i_snitch_regfile.mem\[230\]
+ net3107 i_snitch.i_snitch_regfile.mem\[134\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y
+ i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B
+ VPWR VGND sg13g2_nor2_1
XFILLER_14_802 VPWR VGND sg13g2_fill_1
XFILLER_25_150 VPWR VGND sg13g2_decap_8
XFILLER_26_684 VPWR VGND sg13g2_decap_8
Xheichips25_snitch_wrapper_29 VPWR VGND uio_oe[3] sg13g2_tiehi
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2702 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X
+ VPWR i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C
+ VGND i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y
+ sg13g2_o21ai_1
Xdata_pdata\[20\]_sg13g2_dfrbpq_1_Q net3233 VGND VPWR data_pdata\[20\]_sg13g2_dfrbpq_1_Q_D
+ data_pdata\[20\] clknet_leaf_23_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[402\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[402\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2467 net2272 net2389 net1164 VPWR VGND sg13g2_a22oi_1
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A_sg13g2_nor2_1_Y
+ net3147 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_96_838 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[43\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[267\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
XFILLER_95_326 VPWR VGND sg13g2_decap_4
XFILLER_1_783 VPWR VGND sg13g2_decap_8
XFILLER_76_551 VPWR VGND sg13g2_fill_2
XFILLER_48_242 VPWR VGND sg13g2_fill_1
XFILLER_64_746 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_44_492 VPWR VGND sg13g2_fill_2
XFILLER_20_816 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[126\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[126\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_32_676 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[225\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[225\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net444 net2331 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[276\]_sg13g2_dfrbpq_1_Q_D VGND net2261 net2321
+ sg13g2_o21ai_1
XFILLER_75_2 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[73\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[73\]
+ i_snitch.i_snitch_regfile.mem\[105\] net3123 i_snitch.i_snitch_regfile.mem\[73\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_120_clk clknet_5_4__leaf_clk clknet_leaf_120_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2
+ VGND net2572 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xshift_reg_q\[25\]_sg13g2_dfrbpq_1_Q net3187 VGND VPWR net516 shift_reg_q\[25\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
XFILLER_28_1025 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[215\]_sg13g2_dfrbpq_1_Q_D VGND net2249 net2335
+ sg13g2_o21ai_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[273\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_xnor2_1
XFILLER_100_147 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[144\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_39_220 VPWR VGND sg13g2_fill_2
XFILLER_95_882 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_inv_1_A
+ i_req_register.data_o\[39\]_sg13g2_o21ai_1_Y_A2 net1149 VPWR VGND sg13g2_inv_2
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net456 net2319 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[50\] VGND sg13g2_inv_1
XFILLER_28_949 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ net2748 i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
XFILLER_54_223 VPWR VGND sg13g2_fill_2
XFILLER_27_437 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[494\]_sg13g2_o21ai_1_A1 net2964 VPWR i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[494\] net2804 sg13g2_o21ai_1
XFILLER_54_267 VPWR VGND sg13g2_fill_1
XFILLER_36_960 VPWR VGND sg13g2_fill_1
XFILLER_42_418 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2419 i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[18\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_23_610 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[422\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[422\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2381 net1101 net2899 net2862 VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2599 i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[14\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.inst_addr_o\[14\] net2527 VPWR VGND sg13g2_xnor2_1
XFILLER_50_451 VPWR VGND sg13g2_decap_4
XFILLER_11_816 VPWR VGND sg13g2_fill_2
XFILLER_22_142 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y
+ VGND VPWR net2543 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_a21oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[22\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net3174 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[283\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[283\] VGND sg13g2_inv_1
Xclkbuf_leaf_111_clk clknet_5_5__leaf_clk clknet_leaf_111_clk VPWR VGND sg13g2_buf_8
XFILLER_105_910 VPWR VGND sg13g2_decap_8
Xfanout3229 net3249 net3229 VPWR VGND sg13g2_buf_8
Xfanout3207 net3211 net3207 VPWR VGND sg13g2_buf_8
Xfanout3218 net3225 net3218 VPWR VGND sg13g2_buf_8
XFILLER_104_420 VPWR VGND sg13g2_decap_8
XFILLER_81_1005 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ net1154 VGND sg13g2_inv_1
Xfanout2517 net2518 net2517 VPWR VGND sg13g2_buf_8
Xfanout2506 net2507 net2506 VPWR VGND sg13g2_buf_8
XFILLER_105_987 VPWR VGND sg13g2_decap_8
XFILLER_104_442 VPWR VGND sg13g2_fill_2
Xfanout2539 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y
+ net2539 VPWR VGND sg13g2_buf_8
XFILLER_89_153 VPWR VGND sg13g2_decap_8
XFILLER_78_827 VPWR VGND sg13g2_fill_1
Xfanout2528 net2529 net2528 VPWR VGND sg13g2_buf_8
Xhold393 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net425 sg13g2_dlygate4sd3_1
XFILLER_77_337 VPWR VGND sg13g2_fill_2
XFILLER_86_860 VPWR VGND sg13g2_decap_8
XFILLER_100_681 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y
+ VGND VPWR net2516 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[39\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2427 sg13g2_a21oi_1
XFILLER_46_702 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[313\]_sg13g2_o21ai_1_A1 net2935 VPWR i_snitch.i_snitch_regfile.mem\[313\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[313\] net2810 sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[146\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[146\] clknet_leaf_91_clk sg13g2_dfrbpq_1
Xhold1060 i_snitch.i_snitch_regfile.mem\[218\] VPWR VGND net1092 sg13g2_dlygate4sd3_1
XFILLER_19_938 VPWR VGND sg13g2_decap_8
XFILLER_100_692 VPWR VGND sg13g2_fill_1
XFILLER_73_554 VPWR VGND sg13g2_fill_1
XFILLER_73_532 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1
+ i_snitch.i_snitch_regfile.mem\[57\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y VPWR
+ i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[281\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X sg13g2_o21ai_1
Xhold1082 i_snitch.i_snitch_regfile.mem\[263\] VPWR VGND net1114 sg13g2_dlygate4sd3_1
Xhold1093 i_snitch.i_snitch_regfile.mem\[382\] VPWR VGND net1125 sg13g2_dlygate4sd3_1
XFILLER_34_908 VPWR VGND sg13g2_fill_1
Xhold1071 i_snitch.i_snitch_regfile.mem\[70\] VPWR VGND net1103 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1 net3020 i_snitch.i_snitch_regfile.mem\[401\]
+ i_snitch.i_snitch_regfile.mem\[433\] i_snitch.i_snitch_regfile.mem\[465\] i_snitch.i_snitch_regfile.mem\[497\]
+ net2992 i_snitch.i_snitch_regfile.mem\[401\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
XFILLER_45_278 VPWR VGND sg13g2_decap_8
XFILLER_33_407 VPWR VGND sg13g2_decap_4
XFILLER_73_598 VPWR VGND sg13g2_fill_1
XFILLER_61_749 VPWR VGND sg13g2_decap_4
Xi_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y i_snitch.gpr_waddr\[6\]
+ data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y i_snitch.gpr_waddr\[7\] i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
XFILLER_45_289 VPWR VGND sg13g2_fill_2
XFILLER_26_470 VPWR VGND sg13g2_decap_4
XFILLER_42_985 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[23\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y
+ i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
XFILLER_9_135 VPWR VGND sg13g2_decap_4
Xrebuffer5 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ net37 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C net2312 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2
+ i_req_arb.data_i\[44\] i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
XFILLER_10_871 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2603 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_102_clk clknet_5_19__leaf_clk clknet_leaf_102_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N VPWR VGND sg13g2_nor3_1
XFILLER_69_805 VPWR VGND sg13g2_decap_4
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_68_337 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[351\]_sg13g2_dfrbpq_1_Q_D VGND net2242 net2400
+ sg13g2_o21ai_1
XFILLER_1_580 VPWR VGND sg13g2_decap_8
XFILLER_84_819 VPWR VGND sg13g2_fill_2
XFILLER_84_808 VPWR VGND sg13g2_fill_1
XFILLER_3_98 VPWR VGND sg13g2_decap_8
XFILLER_83_307 VPWR VGND sg13g2_fill_2
XFILLER_92_885 VPWR VGND sg13g2_decap_8
XFILLER_91_362 VPWR VGND sg13g2_fill_1
XFILLER_64_554 VPWR VGND sg13g2_fill_2
XFILLER_24_407 VPWR VGND sg13g2_fill_2
XFILLER_17_470 VPWR VGND sg13g2_fill_2
XFILLER_51_259 VPWR VGND sg13g2_fill_1
XFILLER_51_248 VPWR VGND sg13g2_decap_8
XFILLER_80_0 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A i_snitch.i_snitch_regfile.mem\[113\]
+ net2997 i_snitch.i_snitch_regfile.mem\[113\]_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
XFILLER_105_217 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[166\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[166\] clknet_leaf_86_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_nand2b_1_A_N_Y
+ net121 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\] VPWR
+ VGND sg13g2_nand2b_1
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2
+ i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y net3088
+ i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y i_snitch.i_snitch_regfile.mem\[412\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X
+ net2795 net2912 i_snitch.i_snitch_regfile.mem\[322\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ VPWR VGND sg13g2_and2_1
Xi_snitch.i_snitch_regfile.mem\[263\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2 VGND VPWR
+ net2935 i_snitch.i_snitch_regfile.mem\[263\]_sg13g2_mux4_1_A0_X i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y sg13g2_a21oi_1
XFILLER_102_968 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_D
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A
+ net2744 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_nor4_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y
+ VGND VPWR net3082 net100 i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A
+ i_req_arb.data_i\[43\] sg13g2_a21oi_1
XFILLER_86_167 VPWR VGND sg13g2_fill_1
XFILLER_68_893 VPWR VGND sg13g2_fill_1
XFILLER_83_830 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VGND net2425 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_27_256 VPWR VGND sg13g2_decap_8
XFILLER_103_77 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N_sg13g2_nand3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[6\]_sg13g2_mux2_1_A1_X
+ net2926 net3036 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand3_1
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ net48 i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y
+ i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y
+ VGND VPWR net34 sg13g2_nor4_2
Xrsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[26\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1330 net3067 net1169 VPWR VGND sg13g2_a22oi_1
XFILLER_70_546 VPWR VGND sg13g2_fill_1
XFILLER_70_535 VPWR VGND sg13g2_decap_8
XFILLER_55_587 VPWR VGND sg13g2_fill_1
XFILLER_43_749 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[485\]_sg13g2_nor3_1_A net1249 net2854 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[485\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_50_292 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A VGND
+ VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A_X
+ net2496 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X sg13g2_or2_1
Xi_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[213\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2789
+ net2669 VPWR VGND sg13g2_nand2_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[256\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X i_snitch.i_snitch_regfile.mem\[384\]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ sg13g2_a221oi_1
Xfanout3004 net3006 net3004 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[462\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[462\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2373 net1096 net2687 net2741 VPWR VGND sg13g2_a22oi_1
Xfanout3037 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_Y
+ net3037 VPWR VGND sg13g2_buf_2
Xfanout3026 net3027 net3026 VPWR VGND sg13g2_buf_8
Xfanout3015 net3025 net3015 VPWR VGND sg13g2_buf_8
Xfanout3059 net3062 net3059 VPWR VGND sg13g2_buf_8
Xfanout2303 net2304 net2303 VPWR VGND sg13g2_buf_8
Xfanout2325 net2326 net2325 VPWR VGND sg13g2_buf_8
Xfanout2314 net2315 net2314 VPWR VGND sg13g2_buf_8
XFILLER_3_878 VPWR VGND sg13g2_decap_8
XFILLER_2_355 VPWR VGND sg13g2_fill_2
Xfanout3048 net3049 net3048 VPWR VGND sg13g2_buf_8
XFILLER_105_784 VPWR VGND sg13g2_decap_8
Xfanout2336 net2339 net2336 VPWR VGND sg13g2_buf_8
Xfanout2358 i_snitch.sb_d\[2\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y
+ net2358 VPWR VGND sg13g2_buf_8
Xfanout2347 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2347 VPWR VGND sg13g2_buf_8
Xfanout2369 net2371 net2369 VPWR VGND sg13g2_buf_8
XFILLER_104_294 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.pc_d\[18\]_sg13g2_mux2_1_A1 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1 i_snitch.pc_d\[18\]
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_A1 i_snitch.pc_d\[18\]_sg13g2_mux2_1_A1_X VPWR
+ VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[317\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2779
+ net2654 VPWR VGND sg13g2_nand2_1
XFILLER_77_167 VPWR VGND sg13g2_fill_2
XFILLER_93_649 VPWR VGND sg13g2_decap_4
XFILLER_74_852 VPWR VGND sg13g2_fill_1
XFILLER_74_841 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VGND i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ net230 sg13g2_o21ai_1
XFILLER_73_362 VPWR VGND sg13g2_fill_1
XFILLER_46_587 VPWR VGND sg13g2_fill_1
XFILLER_18_278 VPWR VGND sg13g2_fill_2
XFILLER_34_727 VPWR VGND sg13g2_fill_2
Xshift_reg_q\[8\]_sg13g2_nor2_1_A net503 net2735 shift_reg_q\[8\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_61_568 VPWR VGND sg13g2_decap_4
XFILLER_14_440 VPWR VGND sg13g2_fill_1
XFILLER_33_237 VPWR VGND sg13g2_decap_4
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[27\] net1065 net2915 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[27\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1 net3005 i_snitch.i_snitch_regfile.mem\[405\]
+ i_snitch.i_snitch_regfile.mem\[437\] i_snitch.i_snitch_regfile.mem\[469\] i_snitch.i_snitch_regfile.mem\[501\]
+ net2978 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[186\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[186\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[353\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[353\]
+ net2951 sg13g2_o21ai_1
XFILLER_41_281 VPWR VGND sg13g2_fill_1
XFILLER_42_793 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2 i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1 i_snitch.inst_addr_o\[29\] i_snitch.pc_d\[26\]_sg13g2_a21oi_1_Y_B1
+ i_snitch.inst_addr_o\[26\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1
+ VPWR i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_Y
+ VGND i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C
+ sg13g2_o21ai_1
XFILLER_5_182 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_dfrbpq_1_Q net3224 VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[34\] clknet_leaf_109_clk sg13g2_dfrbpq_1
XFILLER_97_922 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y
+ net2565 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A
+ VPWR VGND sg13g2_nor2_1
XFILLER_69_624 VPWR VGND sg13g2_fill_2
Xfanout2881 net2883 net2881 VPWR VGND sg13g2_buf_8
Xfanout2870 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X net2870
+ VPWR VGND sg13g2_buf_8
XFILLER_97_999 VPWR VGND sg13g2_decap_8
Xfanout2892 net2896 net2892 VPWR VGND sg13g2_buf_8
XFILLER_49_392 VPWR VGND sg13g2_fill_1
XFILLER_65_885 VPWR VGND sg13g2_fill_2
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2
+ VPWR VGND sg13g2_nor2b_1
Xstrb_reg_q\[4\]_sg13g2_dfrbpq_1_Q net3189 VGND VPWR net473 strb_reg_q\[4\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
XFILLER_20_432 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1
+ VGND i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[348\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2655 VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2560 i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1
+ net2720 net3074 i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X
+ VGND VPWR i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1
+ i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B
+ net2717 sg13g2_or2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q
+ net3203 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[24\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
XFILLER_106_548 VPWR VGND sg13g2_fill_1
XFILLER_106_537 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X
+ net2562 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_and2_1
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_102_765 VPWR VGND sg13g2_fill_1
XFILLER_101_231 VPWR VGND sg13g2_decap_8
XFILLER_88_966 VPWR VGND sg13g2_decap_8
XFILLER_102_776 VPWR VGND sg13g2_fill_1
XFILLER_59_178 VPWR VGND sg13g2_fill_2
Xdata_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[373\]_sg13g2_o21ai_1_A1 net2969 VPWR i_snitch.i_snitch_regfile.mem\[373\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[373\] net2802 sg13g2_o21ai_1
XFILLER_28_510 VPWR VGND sg13g2_decap_8
XFILLER_71_800 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2 VGND VPWR
+ net2934 i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[52\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[148\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y sg13g2_a21oi_1
XFILLER_55_351 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2854
+ net2661 VPWR VGND sg13g2_nand2_1
XFILLER_70_321 VPWR VGND sg13g2_fill_2
XFILLER_16_727 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A_Y net2950 i_snitch.i_snitch_regfile.mem\[70\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ net2942 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2
+ net2632 VPWR i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VGND net2635 i_snitch.i_snitch_regfile.mem\[269\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_15_248 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[301\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[301\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2689 net2779 net2317 net1260 VPWR VGND sg13g2_a22oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[11\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q net3320 VGND VPWR i_snitch.i_snitch_regfile.mem\[54\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[54\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_12_988 VPWR VGND sg13g2_fill_1
XFILLER_87_1000 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[275\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2891
+ net2673 VPWR VGND sg13g2_nand2_1
XFILLER_99_77 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[508\]_sg13g2_o21ai_1_A1 net2963 VPWR i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[508\] net2801 sg13g2_o21ai_1
XFILLER_97_207 VPWR VGND sg13g2_decap_4
XFILLER_79_900 VPWR VGND sg13g2_fill_1
XFILLER_3_653 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_79_944 VPWR VGND sg13g2_decap_8
XFILLER_2_141 VPWR VGND sg13g2_fill_1
XFILLER_94_903 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_78_476 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1 VPWR VGND
+ i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_a21oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[297\]_sg13g2_o21ai_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[329\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y net2919
+ sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[379\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2878
+ net2658 VPWR VGND sg13g2_nand2_1
XFILLER_94_1015 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[27\]_sg13g2_a21oi_1_Y_A1
+ net2303 i_snitch.pc_d\[27\] net57 sg13g2_a21oi_1
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_34_546 VPWR VGND sg13g2_fill_1
XFILLER_61_387 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q
+ net3253 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[44\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
XFILLER_21_218 VPWR VGND sg13g2_fill_2
XFILLER_22_719 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y
+ VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[8\]_sg13g2_mux2_1_A1_1_X
+ net2535 i_snitch.pc_d\[1\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B
+ i_snitch.inst_addr_o\[1\] sg13g2_a21oi_1
XFILLER_9_42 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[395\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y
+ VPWR VGND sg13g2_and3_1
Xhold904 i_snitch.i_snitch_regfile.mem\[428\] VPWR VGND net936 sg13g2_dlygate4sd3_1
Xhold937 i_snitch.i_snitch_regfile.mem\[500\] VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold926 i_snitch.i_snitch_regfile.mem\[253\] VPWR VGND net958 sg13g2_dlygate4sd3_1
Xhold915 i_snitch.i_snitch_regfile.mem\[334\] VPWR VGND net947 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B
+ net2576 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_2
Xhold959 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] VPWR
+ VGND net991 sg13g2_dlygate4sd3_1
Xhold948 i_snitch.i_snitch_regfile.mem\[208\] VPWR VGND net980 sg13g2_dlygate4sd3_1
XFILLER_103_518 VPWR VGND sg13g2_fill_2
XFILLER_88_229 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1 net3004 i_snitch.i_snitch_regfile.mem\[409\]
+ i_snitch.i_snitch_regfile.mem\[441\] i_snitch.i_snitch_regfile.mem\[473\] i_snitch.i_snitch_regfile.mem\[505\]
+ net2977 i_snitch.i_snitch_regfile.mem\[409\]_sg13g2_mux4_1_A0_1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[306\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[306\] VGND sg13g2_inv_1
XFILLER_85_969 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q net3270 VGND VPWR i_snitch.i_snitch_regfile.mem\[74\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[74\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_91_clk clknet_5_20__leaf_clk clknet_leaf_91_clk VPWR VGND sg13g2_buf_8
XFILLER_100_56 VPWR VGND sg13g2_decap_8
XFILLER_60_27 VPWR VGND sg13g2_fill_1
Xdata_pdata\[6\]_sg13g2_mux2_1_A1 rsp_data_q\[6\] net719 net3051 data_pdata\[6\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2819 i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
Xshift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y VGND VPWR net2728 shift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2
+ shift_reg_q\[25\]_sg13g2_dfrbpq_1_Q_D shift_reg_q\[25\]_sg13g2_nor2_1_A_Y sg13g2_a21oi_1
XFILLER_21_785 VPWR VGND sg13g2_decap_4
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2297 net1169 net2495 net1274 VPWR VGND sg13g2_a22oi_1
XFILLER_5_907 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[467\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[93\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[125\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
XFILLER_106_301 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2604 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y
+ VGND VPWR i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_106_378 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[357\]_sg13g2_nor3_1_A net1337 net2878 i_snitch.sb_d\[11\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B
+ net3087 net2719 i_req_arb.data_i\[40\] VPWR VGND sg13g2_a22oi_1
XFILLER_0_667 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2 i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0_X
+ net2936 net2930 i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_87_284 VPWR VGND sg13g2_decap_8
XFILLER_48_649 VPWR VGND sg13g2_fill_2
XFILLER_56_660 VPWR VGND sg13g2_decap_4
XFILLER_47_159 VPWR VGND sg13g2_decap_8
XFILLER_18_40 VPWR VGND sg13g2_fill_2
XFILLER_28_340 VPWR VGND sg13g2_fill_2
XFILLER_28_351 VPWR VGND sg13g2_fill_1
XFILLER_29_852 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2558 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_mux2_1_A1
+ net775 net608 net2239 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_82_clk clknet_5_29__leaf_clk clknet_leaf_82_clk VPWR VGND sg13g2_buf_8
Xrsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ net1294 VGND sg13g2_inv_1
Xi_req_arb.data_i\[44\]_sg13g2_a21o_1_B1 net100 net3080 i_req_arb.data_i\[44\] i_req_arb.data_i\[44\]_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_1
XFILLER_54_1021 VPWR VGND sg13g2_decap_8
Xuio_out_sg13g2_buf_1_X_3 i_req_register.data_o\[45\] net16 VPWR VGND sg13g2_buf_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A
+ net2483 i_snitch.i_snitch_regfile.mem\[286\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net2746 i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_7_222 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[149\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[61\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2768
+ net2654 VPWR VGND sg13g2_nand2_1
XFILLER_50_60 VPWR VGND sg13g2_fill_2
XFILLER_8_778 VPWR VGND sg13g2_fill_1
XFILLER_7_266 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2 i_snitch.inst_addr_o\[20\]
+ VPWR i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2_Y VGND net2305 i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1
+ sg13g2_o21ai_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_nand2_1
XFILLER_7_277 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[341\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[341\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2401 net948 net2472 net2269 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1_sg13g2_inv_1_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[45\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1
+ net1074 VGND sg13g2_inv_1
XFILLER_4_962 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q net3285 VGND VPWR i_snitch.i_snitch_regfile.mem\[94\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[94\] clknet_leaf_87_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\] net620 net2617
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2286
+ net2467 VPWR VGND sg13g2_nand2_1
XFILLER_79_774 VPWR VGND sg13g2_fill_2
XFILLER_94_755 VPWR VGND sg13g2_fill_1
XFILLER_94_722 VPWR VGND sg13g2_fill_1
XFILLER_66_413 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1
+ net2501 VGND sg13g2_inv_1
XFILLER_19_373 VPWR VGND sg13g2_decap_4
XFILLER_19_384 VPWR VGND sg13g2_fill_1
Xi_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y VPWR VGND net2934
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 i_snitch.i_snitch_regfile.mem\[50\]_sg13g2_a22oi_1_A1_Y
+ net3088 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2 i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_or3_1_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1
+ VPWR VGND sg13g2_or3_1
XFILLER_46_192 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_73_clk clknet_5_25__leaf_clk clknet_leaf_73_clk VPWR VGND sg13g2_buf_8
XFILLER_90_994 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[0\]_sg13g2_dfrbpq_1_Q net3230 VGND VPWR rsp_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[0\] clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_22_505 VPWR VGND sg13g2_fill_2
XFILLER_34_387 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[494\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2275
+ net2459 VPWR VGND sg13g2_nand2_1
Xdata_pdata\[18\]_sg13g2_mux2_1_A0 data_pdata\[18\] data_pdata\[26\] net3156 data_pdata\[18\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold701 i_snitch.i_snitch_regfile.mem\[329\] VPWR VGND net733 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_or2_1_A_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xhold712 i_snitch.i_snitch_regfile.mem\[463\] VPWR VGND net744 sg13g2_dlygate4sd3_1
Xhold745 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\] VPWR
+ VGND net777 sg13g2_dlygate4sd3_1
Xhold734 i_snitch.i_snitch_regfile.mem\[88\] VPWR VGND net766 sg13g2_dlygate4sd3_1
Xhold723 data_pdata\[19\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net755 sg13g2_dlygate4sd3_1
XFILLER_104_816 VPWR VGND sg13g2_decap_8
XFILLER_103_315 VPWR VGND sg13g2_decap_8
Xhold778 data_pdata\[16\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net810 sg13g2_dlygate4sd3_1
Xhold767 data_pdata\[22\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net799 sg13g2_dlygate4sd3_1
Xhold756 i_snitch.i_snitch_regfile.mem\[457\] VPWR VGND net788 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1
+ net2725 i_snitch.inst_addr_o\[16\] i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
Xhold789 i_snitch.i_snitch_regfile.mem\[40\] VPWR VGND net821 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_nand2b_1_B i_snitch.i_snitch_lsu.metadata_q\[1\]_sg13g2_nand2b_1_B_Y
+ i_snitch.i_snitch_lsu.metadata_q\[1\] net3151 VPWR VGND sg13g2_nand2b_1
XFILLER_97_593 VPWR VGND sg13g2_decap_8
XFILLER_58_958 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]_sg13g2_dfrbpq_1_Q
+ net3186 VGND VPWR net572 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[11\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2778 i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2908 net2430 i_snitch.i_snitch_regfile.mem\[292\]_sg13g2_dfrbpq_1_Q_D net2476
+ sg13g2_a221oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\] net577 net2623
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[10\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[92\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2784
+ net2656 VPWR VGND sg13g2_nand2_1
XFILLER_84_287 VPWR VGND sg13g2_decap_8
XFILLER_44_107 VPWR VGND sg13g2_decap_4
XFILLER_26_822 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2586 i_snitch.pc_d\[11\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2
+ net101 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_64_clk clknet_5_28__leaf_clk clknet_leaf_64_clk VPWR VGND sg13g2_buf_8
XFILLER_53_685 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[361\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[361\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2398 net795 net2686 net2880 VPWR VGND sg13g2_a22oi_1
XFILLER_38_1016 VPWR VGND sg13g2_decap_8
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2722 i_snitch.inst_addr_o\[11\] sg13g2_a21oi_2
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q net3250 VGND VPWR i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_lsu.metadata_q\[0\] clknet_leaf_15_clk sg13g2_dfrbpq_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y
+ net2501 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ net2508 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_2
Xi_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[405\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ net2723 i_snitch.inst_addr_o\[21\] sg13g2_a21oi_2
Xi_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[285\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[21\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2596 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_nand2_1
XFILLER_84_1003 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
XFILLER_106_175 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1
+ net88 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y
+ net2565 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[362\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[362\]
+ net3132 i_snitch.i_snitch_regfile.mem\[362\]_sg13g2_a21oi_1_A1_Y net2942 sg13g2_a21oi_1
XFILLER_96_56 VPWR VGND sg13g2_decap_8
XFILLER_88_571 VPWR VGND sg13g2_decap_4
XFILLER_76_711 VPWR VGND sg13g2_decap_8
XFILLER_1_965 VPWR VGND sg13g2_decap_8
XFILLER_103_893 VPWR VGND sg13g2_decap_8
XFILLER_49_958 VPWR VGND sg13g2_fill_2
XFILLER_0_475 VPWR VGND sg13g2_decap_8
XFILLER_102_392 VPWR VGND sg13g2_decap_8
XFILLER_76_755 VPWR VGND sg13g2_fill_1
XFILLER_64_917 VPWR VGND sg13g2_fill_1
XFILLER_57_980 VPWR VGND sg13g2_fill_1
XFILLER_17_800 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y
+ net2552 VPWR i_snitch.pc_d\[24\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1
+ VGND net2745 i_snitch.i_snitch_regfile.mem\[152\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
Xclkbuf_leaf_55_clk clknet_5_30__leaf_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2361 net1013 net2900 net2768 VPWR VGND sg13g2_a22oi_1
Xrsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[24\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1167 net3063 net907 VPWR VGND sg13g2_a22oi_1
XFILLER_16_343 VPWR VGND sg13g2_fill_1
XFILLER_17_877 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[141\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A
+ net73 net2724 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[489\]_sg13g2_dfrbpq_1_Q_D VGND net2299 net2366
+ sg13g2_o21ai_1
XFILLER_31_368 VPWR VGND sg13g2_fill_2
XFILLER_84_7 VPWR VGND sg13g2_fill_2
XFILLER_6_21 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[39\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[39\]
+ net2824 i_snitch.i_snitch_regfile.mem\[39\]_sg13g2_a21oi_1_A1_Y net2821 sg13g2_a21oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_dfrbpq_1_Q
+ net3187 VGND VPWR net638 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
XFILLER_99_825 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_6_98 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nand2b_1_A_N i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_nand2b_1_A_N_Y
+ net3026 i_snitch.i_snitch_regfile.mem\[67\] VPWR VGND sg13g2_nand2b_1
Xi_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[428\]_sg13g2_dfrbpq_1_Q_D VGND net2277 net2379
+ sg13g2_o21ai_1
XFILLER_101_819 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[381\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[381\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2395 net1022 net2470 net2250 VPWR VGND sg13g2_a22oi_1
XFILLER_66_232 VPWR VGND sg13g2_fill_2
XFILLER_66_221 VPWR VGND sg13g2_decap_8
Xrebuffer26 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A
+ net58 VPWR VGND sg13g2_buf_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X
+ i_snitch.i_snitch_regfile.mem\[51\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y
+ VPWR VGND sg13g2_nor3_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]
+ net3177 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X
+ VPWR VGND sg13g2_mux2_1
Xrebuffer15 i_snitch.i_snitch_regfile.mem\[130\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y
+ net47 VPWR VGND sg13g2_buf_8
Xrebuffer37 i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B
+ net69 VPWR VGND sg13g2_buf_1
Xclkbuf_leaf_46_clk clknet_5_12__leaf_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
Xrebuffer59 i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y net91 VPWR VGND sg13g2_buf_1
Xrebuffer48 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[20\]_sg13g2_mux2_1_A1_X
+ net80 VPWR VGND sg13g2_buf_1
XFILLER_23_836 VPWR VGND sg13g2_decap_8
XFILLER_34_195 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1
+ net2815 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2 VPWR VGND i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp
+ i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y
+ net3172 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[382\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[382\]
+ net3127 i_snitch.i_snitch_regfile.mem\[382\]_sg13g2_a21oi_1_A1_Y net2943 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[34\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2485 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_nor3_1_A_Y net2454 net2765 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_dfrbpq_1_Q_D
+ net2912 sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X
+ i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[388\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y
+ sg13g2_a21oi_1
Xhold520 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[16\] VPWR
+ VGND net552 sg13g2_dlygate4sd3_1
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1
+ net490 i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B VPWR VGND sg13g2_nand2_1
Xhold531 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\] VPWR
+ VGND net563 sg13g2_dlygate4sd3_1
Xhold553 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net585 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[272\]_sg13g2_o21ai_1_A1 net2936 VPWR i_snitch.i_snitch_regfile.mem\[272\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[272\] net2814 sg13g2_o21ai_1
Xhold542 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\] VPWR
+ VGND net574 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[42\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_103_112 VPWR VGND sg13g2_decap_8
Xhold586 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[29\] VPWR
+ VGND net618 sg13g2_dlygate4sd3_1
Xhold597 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[28\] VPWR
+ VGND net629 sg13g2_dlygate4sd3_1
Xhold564 i_snitch.sb_q\[6\] VPWR VGND net596 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[411\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[411\] clknet_leaf_119_clk sg13g2_dfrbpq_1
Xhold575 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net607 sg13g2_dlygate4sd3_1
XFILLER_77_519 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[200\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[200\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2337 net823 net2643 net2791 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2359 net981 net2454 net2255 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[106\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y
+ VGND net2819 i_snitch.i_snitch_regfile.mem\[138\]_sg13g2_mux4_1_A0_X sg13g2_o21ai_1
XFILLER_106_77 VPWR VGND sg13g2_decap_8
XFILLER_103_189 VPWR VGND sg13g2_decap_8
Xhold1231 rsp_data_q\[4\] VPWR VGND net1263 sg13g2_dlygate4sd3_1
Xhold1220 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[34\] VPWR
+ VGND net1252 sg13g2_dlygate4sd3_1
Xhold1242 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[28\] VPWR
+ VGND net1274 sg13g2_dlygate4sd3_1
XFILLER_57_221 VPWR VGND sg13g2_decap_8
XFILLER_46_917 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[9\] net632 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[9\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_100_896 VPWR VGND sg13g2_decap_8
XFILLER_58_799 VPWR VGND sg13g2_fill_2
XFILLER_58_788 VPWR VGND sg13g2_decap_8
Xhold1264 i_snitch.i_snitch_regfile.mem\[437\] VPWR VGND net1296 sg13g2_dlygate4sd3_1
Xhold1253 i_snitch.i_snitch_regfile.mem\[443\] VPWR VGND net1285 sg13g2_dlygate4sd3_1
Xhold1275 i_snitch.i_snitch_regfile.mem\[482\] VPWR VGND net1307 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_37_clk clknet_5_10__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_73_758 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_nand2_1_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_nand2_1_A_Y
+ net426 net2623 VPWR VGND sg13g2_nand2_1
Xhold1286 i_snitch.i_snitch_regfile.mem\[296\] VPWR VGND net1318 sg13g2_dlygate4sd3_1
Xhold1297 i_snitch.i_snitch_regfile.mem\[196\] VPWR VGND net1329 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[337\]_sg13g2_dfrbpq_1_Q_D VGND net2288 net2399
+ sg13g2_o21ai_1
XFILLER_25_173 VPWR VGND sg13g2_decap_4
XFILLER_15_96 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[229\]_sg13g2_nor3_1_A net1368 net2872 i_snitch.sb_d\[7\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[229\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1
+ i_snitch.i_snitch_regfile.mem\[136\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A
+ net86 net2750 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y
+ VPWR VGND sg13g2_nor2b_2
Xi_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1 VGND VPWR i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1_A1
+ net41 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a21o_1_A1_B1 sg13g2_a21oi_1
XFILLER_5_534 VPWR VGND sg13g2_fill_2
Xi_req_arb.data_i\[40\]_sg13g2_inv_1_A i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A net1235
+ VPWR VGND sg13g2_inv_2
XFILLER_1_762 VPWR VGND sg13g2_decap_8
XFILLER_95_316 VPWR VGND sg13g2_decap_4
Xi_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_inv_1_A
+ VPWR i_snitch.i_snitch_regfile.mem\[63\]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[30\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A
+ VGND sg13g2_inv_1
XFILLER_48_232 VPWR VGND sg13g2_decap_4
XFILLER_0_294 VPWR VGND sg13g2_fill_1
Xshift_reg_q\[2\]_sg13g2_dfrbpq_1_Q net3195 VGND VPWR net480 shift_reg_q\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_76_574 VPWR VGND sg13g2_fill_1
XFILLER_37_928 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_28_clk clknet_5_9__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_36_438 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D
+ VPWR VGND sg13g2_or4_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_mux2_1_A1
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\] net647 net2619
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[503\]_sg13g2_dfrbpq_1_Q_D VGND net2248 net2365
+ sg13g2_o21ai_1
XFILLER_20_806 VPWR VGND sg13g2_fill_1
XFILLER_32_688 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q net3294 VGND VPWR i_snitch.i_snitch_regfile.mem\[431\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[431\] clknet_leaf_79_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[60\]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2837 i_snitch.i_snitch_regfile.mem\[156\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1 net3006 i_snitch.i_snitch_regfile.mem\[259\]
+ i_snitch.i_snitch_regfile.mem\[291\] i_snitch.i_snitch_regfile.mem\[323\] i_snitch.i_snitch_regfile.mem\[355\]
+ net2979 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X VPWR VGND sg13g2_mux4_1
Xi_snitch.i_snitch_regfile.mem\[220\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[220\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2336 net970 net2440 net2246 VPWR VGND sg13g2_a22oi_1
XFILLER_9_873 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[78\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[78\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2355 net1091 net2688 net2786 VPWR VGND sg13g2_a22oi_1
XFILLER_99_644 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[246\]_sg13g2_dfrbpq_1_Q_D VGND net2258 net2329
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2408 i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2448 net2866 i_snitch.i_snitch_regfile.mem\[101\]_sg13g2_dfrbpq_1_Q_D net2906
+ sg13g2_a221oi_1
XFILLER_99_688 VPWR VGND sg13g2_decap_8
XFILLER_86_327 VPWR VGND sg13g2_decap_4
XFILLER_100_126 VPWR VGND sg13g2_decap_8
XFILLER_95_861 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A
+ i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[79\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[79\]
+ net2845 i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_a21oi_1_A1_Y net2835 sg13g2_a21oi_1
Xi_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1_sg13g2_nand3_1_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1
+ VPWR VGND sg13g2_nand3_1
XFILLER_28_939 VPWR VGND sg13g2_decap_4
XFILLER_39_276 VPWR VGND sg13g2_decap_8
XFILLER_54_213 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_19_clk clknet_5_6__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_82_577 VPWR VGND sg13g2_decap_8
XFILLER_82_566 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A
+ VPWR VGND sg13g2_nand2b_1
XFILLER_42_408 VPWR VGND sg13g2_decap_4
XFILLER_74_1013 VPWR VGND sg13g2_decap_8
XFILLER_35_471 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[111\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[79\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[111\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[111\]
+ net2952 sg13g2_o21ai_1
XFILLER_23_666 VPWR VGND sg13g2_fill_2
XFILLER_23_688 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2
+ net50 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
XFILLER_10_338 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1
+ net2560 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2_Y
+ VPWR VGND sg13g2_xnor2_1
Xrsp_data_q\[12\]_sg13g2_dfrbpq_1_Q net3240 VGND VPWR rsp_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ rsp_data_q\[12\] clknet_leaf_39_clk sg13g2_dfrbpq_2
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A
+ i_snitch.pc_d\[24\]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X net78 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B
+ VPWR VGND sg13g2_nand3_1
Xfanout3208 net3211 net3208 VPWR VGND sg13g2_buf_2
Xfanout3219 net3220 net3219 VPWR VGND sg13g2_buf_8
Xfanout2518 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X
+ net2518 VPWR VGND sg13g2_buf_8
Xfanout2507 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y
+ net2507 VPWR VGND sg13g2_buf_8
XFILLER_105_966 VPWR VGND sg13g2_decap_8
XFILLER_81_1028 VPWR VGND sg13g2_fill_1
Xfanout2529 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[31\]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A_X
+ net2529 VPWR VGND sg13g2_buf_8
Xhold394 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\] VPWR
+ VGND net426 sg13g2_dlygate4sd3_1
XFILLER_104_498 VPWR VGND sg13g2_fill_1
XFILLER_104_476 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_nor2_1_A net554 net2486 i_snitch.i_snitch_lsu.metadata_q\[0\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_92_319 VPWR VGND sg13g2_decap_8
Xhold1050 i_snitch.i_snitch_regfile.mem\[44\] VPWR VGND net1082 sg13g2_dlygate4sd3_1
Xhold1072 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[13\]
+ VPWR VGND net1104 sg13g2_dlygate4sd3_1
Xhold1061 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] VPWR
+ VGND net1093 sg13g2_dlygate4sd3_1
XFILLER_93_35 VPWR VGND sg13g2_decap_8
Xhold1094 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]
+ VPWR VGND net1126 sg13g2_dlygate4sd3_1
XFILLER_18_427 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q net3274 VGND VPWR i_snitch.i_snitch_regfile.mem\[451\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[451\] clknet_leaf_112_clk sg13g2_dfrbpq_1
Xhold1083 i_snitch.i_snitch_regfile.mem\[77\] VPWR VGND net1115 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[260\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[260\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[240\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[240\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2332 net1058 net2438 net2263 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y
+ net94 net2496 net1380 VPWR VGND sg13g2_a22oi_1
XFILLER_42_964 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_dfrbpq_1_Q_D VGND net2522 net2357
+ sg13g2_o21ai_1
Xrebuffer6 i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y
+ net38 VPWR VGND sg13g2_buf_1
Xi_snitch.i_snitch_regfile.mem\[447\]_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[447\]_sg13g2_o21ai_1_A1_Y VGND i_snitch.i_snitch_regfile.mem\[447\]
+ net2812 sg13g2_o21ai_1
XFILLER_6_887 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]_sg13g2_dfrbpq_1_Q
+ net3240 VGND VPWR net1062 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[25\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_96_614 VPWR VGND sg13g2_fill_2
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y
+ VGND VPWR net2420 i_snitch.i_snitch_regfile.mem\[304\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
XFILLER_68_349 VPWR VGND sg13g2_decap_4
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_97_1013 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2
+ i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A i_snitch.pc_d\[20\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[10\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2482 i_snitch.i_snitch_regfile.mem\[308\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2532 VPWR VGND sg13g2_a22oi_1
XFILLER_92_864 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A i_snitch.pc_d\[15\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y
+ i_snitch.pc_d\[16\]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y VPWR VGND sg13g2_and3_1
XFILLER_36_246 VPWR VGND sg13g2_decap_8
XFILLER_64_588 VPWR VGND sg13g2_decap_8
XFILLER_73_0 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[132\]_sg13g2_nor3_1_A net1247 net2890 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[132\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 VPWR
+ VGND sg13g2_nor3_1
Xstrb_reg_q\[6\]_sg13g2_nor2_1_A net442 net2729 strb_reg_q\[6\]_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nor2_1
XFILLER_8_191 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_8_clk clknet_5_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_B1
+ net893 net2310 VPWR VGND sg13g2_nand2_1
XFILLER_99_463 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q net3318 VGND VPWR i_snitch.i_snitch_regfile.mem\[471\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[471\] clknet_leaf_67_clk sg13g2_dfrbpq_1
XFILLER_102_947 VPWR VGND sg13g2_decap_8
Xdata_pdata\[14\]_sg13g2_nand2b_1_B data_pdata\[14\]_sg13g2_nand2b_1_B_Y data_pdata\[14\]
+ net3162 VPWR VGND sg13g2_nand2b_1
XFILLER_87_669 VPWR VGND sg13g2_fill_2
XFILLER_47_28 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[390\] VGND sg13g2_inv_1
XFILLER_55_544 VPWR VGND sg13g2_fill_2
XFILLER_103_56 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2
+ net2580 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_a21o_1
XFILLER_83_886 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[510\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[510\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net453 net2369 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A_Y net2841 i_snitch.i_snitch_regfile.mem\[476\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[508\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_42_249 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2 i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y
+ VGND net2839 i_snitch.i_snitch_regfile.mem\[151\]_sg13g2_mux4_1_A0_1_X sg13g2_o21ai_1
XFILLER_11_614 VPWR VGND sg13g2_fill_2
Xdata_pdata\[13\]_sg13g2_dfrbpq_1_Q net3202 VGND VPWR net726 data_pdata\[13\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C_sg13g2_and3_1_X
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C
+ net3076 net3079 i_snitch.i_snitch_regfile.mem\[34\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_and3_1
Xi_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1 i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[399\]_sg13g2_mux4_1_A0_X net3097 i_snitch.i_snitch_regfile.mem\[303\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[335\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y VPWR VGND
+ sg13g2_a22oi_1
Xfanout3005 net3006 net3005 VPWR VGND sg13g2_buf_8
Xfanout3016 net3018 net3016 VPWR VGND sg13g2_buf_8
Xfanout3027 net3032 net3027 VPWR VGND sg13g2_buf_8
XFILLER_105_763 VPWR VGND sg13g2_decap_8
Xfanout2304 net106 net2304 VPWR VGND sg13g2_buf_8
Xi_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0 net3136 i_snitch.i_snitch_regfile.mem\[145\]
+ i_snitch.i_snitch_regfile.mem\[177\] i_snitch.i_snitch_regfile.mem\[209\] i_snitch.i_snitch_regfile.mem\[241\]
+ net3112 i_snitch.i_snitch_regfile.mem\[145\]_sg13g2_mux4_1_A0_X VPWR VGND sg13g2_mux4_1
Xfanout2326 net2327 net2326 VPWR VGND sg13g2_buf_8
Xfanout2315 i_snitch.sb_d\[9\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2315 VPWR VGND sg13g2_buf_8
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xfanout3038 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y net3038 VPWR VGND sg13g2_buf_8
Xfanout3049 net3052 net3049 VPWR VGND sg13g2_buf_8
XFILLER_104_273 VPWR VGND sg13g2_decap_8
XFILLER_78_614 VPWR VGND sg13g2_decap_8
Xfanout2348 i_snitch.sb_d\[4\]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y
+ net2348 VPWR VGND sg13g2_buf_8
Xfanout2359 net2360 net2359 VPWR VGND sg13g2_buf_8
Xfanout2337 net2338 net2337 VPWR VGND sg13g2_buf_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X
+ rsp_data_q\[22\] net1126 net2913 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[22\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
XFILLER_93_639 VPWR VGND sg13g2_fill_2
XFILLER_101_980 VPWR VGND sg13g2_decap_8
XFILLER_19_725 VPWR VGND sg13g2_decap_8
XFILLER_61_503 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q net3323 VGND VPWR i_snitch.i_snitch_regfile.mem\[119\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[119\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_42_750 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y
+ net2628 i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.pc_d\[3\]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y
+ net2756 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[279\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[279\] VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q net3321 VGND VPWR i_snitch.i_snitch_regfile.mem\[491\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[491\] clknet_leaf_64_clk sg13g2_dfrbpq_1
Xi_req_arb.data_i\[38\]_sg13g2_dfrbpq_1_Q net3261 VGND VPWR i_snitch.pc_d\[3\] i_req_arb.data_i\[38\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
Xi_snitch.i_snitch_regfile.mem\[280\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[280\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2325 net1118 net2666 net2893 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y
+ VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_inv_1_A_Y
+ net2617 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[193\]_sg13g2_nand2_1_A i_snitch.i_snitch_regfile.mem\[193\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A
+ net452 net2337 VPWR VGND sg13g2_nand2_1
Xshift_reg_q\[18\]_sg13g2_dfrbpq_1_Q net3199 VGND VPWR net509 shift_reg_q\[18\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_97_901 VPWR VGND sg13g2_decap_8
XFILLER_96_422 VPWR VGND sg13g2_decap_4
XFILLER_96_400 VPWR VGND sg13g2_fill_2
XFILLER_69_614 VPWR VGND sg13g2_fill_2
XFILLER_97_978 VPWR VGND sg13g2_decap_8
Xfanout2882 net2883 net2882 VPWR VGND sg13g2_buf_8
Xfanout2860 net2861 net2860 VPWR VGND sg13g2_buf_8
Xfanout2871 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X net2871
+ VPWR VGND sg13g2_buf_8
XFILLER_84_617 VPWR VGND sg13g2_decap_8
XFILLER_68_179 VPWR VGND sg13g2_fill_2
XFILLER_68_168 VPWR VGND sg13g2_fill_1
Xfanout2893 net2894 net2893 VPWR VGND sg13g2_buf_8
XFILLER_77_691 VPWR VGND sg13g2_fill_2
XFILLER_64_341 VPWR VGND sg13g2_fill_1
XFILLER_80_845 VPWR VGND sg13g2_fill_2
XFILLER_80_834 VPWR VGND sg13g2_fill_2
XFILLER_80_823 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1 VPWR VGND i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C_Y i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1
+ i_req_arb.data_i\[43\] i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_Y
+ i_snitch.pc_d\[8\]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A_X sg13g2_a221oi_1
Xi_snitch.i_snitch_regfile.mem\[84\]_sg13g2_mux2_1_A0 i_snitch.i_snitch_regfile.mem\[84\]
+ i_snitch.i_snitch_regfile.mem\[116\] net3138 i_snitch.i_snitch_regfile.mem\[84\]_sg13g2_mux2_1_A0_X
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[415\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_a22oi_1_B2_Y
+ net2388 net597 net2646 net3039 VPWR VGND sg13g2_a22oi_1
XFILLER_37_588 VPWR VGND sg13g2_decap_4
XFILLER_52_569 VPWR VGND sg13g2_fill_2
XFILLER_24_249 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ net2712 i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y
+ VGND VPWR net2551 i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[19\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1
+ i_snitch.i_snitch_regfile.mem\[300\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ sg13g2_a21oi_1
XFILLER_80_889 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[22\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net1169 net3063 rsp_data_q\[18\] VPWR VGND sg13g2_a22oi_1
XFILLER_33_750 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q net3314 VGND VPWR i_snitch.i_snitch_regfile.mem\[310\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[310\] clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_106_516 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[416\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[416\]
+ net3010 i_snitch.i_snitch_regfile.mem\[416\]_sg13g2_a21oi_1_A1_Y net2981 sg13g2_a21oi_1
Xi_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1
+ net2709 i_snitch.i_snitch_regfile.mem\[291\]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y
+ VPWR VGND sg13g2_nand2_1
XFILLER_88_945 VPWR VGND sg13g2_decap_8
XFILLER_101_210 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[427\] VGND sg13g2_inv_1
XFILLER_48_809 VPWR VGND sg13g2_fill_2
XFILLER_0_849 VPWR VGND sg13g2_decap_8
XFILLER_75_628 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q net3319 VGND VPWR i_snitch.i_snitch_regfile.mem\[139\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[139\] clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_101_287 VPWR VGND sg13g2_decap_8
XFILLER_68_680 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0
+ VGND net2712 i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y
+ sg13g2_o21ai_1
XFILLER_83_650 VPWR VGND sg13g2_decap_4
XFILLER_74_37 VPWR VGND sg13g2_fill_2
XFILLER_83_683 VPWR VGND sg13g2_fill_1
Xrsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[7\]_sg13g2_dfrbpq_1_Q_D
+ net1300 VGND sg13g2_inv_1
XFILLER_55_374 VPWR VGND sg13g2_fill_2
XFILLER_90_14 VPWR VGND sg13g2_decap_8
XFILLER_70_388 VPWR VGND sg13g2_fill_2
Xdata_pdata\[11\]_sg13g2_mux2_1_A1 rsp_data_q\[11\] net995 net3049 data_pdata\[11\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xshift_reg_q\[6\]_sg13g2_a22oi_1_A1 shift_reg_q\[6\]_sg13g2_a22oi_1_A1_Y i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_mux2_1_A1_1_X
+ net3055 net3045 shift_reg_q\[6\] VPWR VGND sg13g2_a22oi_1
XFILLER_23_271 VPWR VGND sg13g2_fill_1
XFILLER_23_85 VPWR VGND sg13g2_fill_1
Xdata_pdata\[25\]_sg13g2_a21oi_1_A2 VGND VPWR net3155 data_pdata\[25\] data_pdata\[25\]_sg13g2_a21oi_1_A2_Y
+ data_pdata\[17\]_sg13g2_nor2b_1_B_N_Y sg13g2_a21oi_1
XFILLER_99_56 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y
+ i_snitch.i_snitch_regfile.mem\[150\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y
+ net2849 net3096 sg13g2_a21oi_2
XFILLER_3_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[435\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[435\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2463 net2270 net2384 net1255 VPWR VGND sg13g2_a22oi_1
XFILLER_93_414 VPWR VGND sg13g2_decap_8
XFILLER_94_959 VPWR VGND sg13g2_decap_8
XFILLER_93_436 VPWR VGND sg13g2_fill_1
XFILLER_19_522 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D
+ i_req_arb.data_i\[42\]_sg13g2_a221oi_1_A1_Y i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ i_snitch.i_snitch_regfile.mem\[38\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D_Y
+ VPWR VGND i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y
+ sg13g2_nand4_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1
+ net2751 net3084 i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X
+ VPWR VGND sg13g2_a21o_2
XFILLER_74_661 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q net3269 VGND VPWR i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[330\] clknet_leaf_102_clk sg13g2_dfrbpq_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q
+ net3260 VGND VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\]_sg13g2_dfrbpq_1_Q_D
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[12\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
XFILLER_74_672 VPWR VGND sg13g2_fill_1
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_525 VPWR VGND sg13g2_fill_1
XFILLER_62_889 VPWR VGND sg13g2_fill_2
XFILLER_9_21 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ VGND net65 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[436\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[436\]
+ net3023 i_snitch.i_snitch_regfile.mem\[436\]_sg13g2_a21oi_1_A1_Y net2993 sg13g2_a21oi_1
XFILLER_15_794 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[158\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2889
+ net2649 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q net3304 VGND VPWR i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[159\] clknet_leaf_51_clk sg13g2_dfrbpq_1
Xhold905 i_snitch.i_snitch_regfile.mem\[156\] VPWR VGND net937 sg13g2_dlygate4sd3_1
Xhold916 i_snitch.i_snitch_regfile.mem\[341\] VPWR VGND net948 sg13g2_dlygate4sd3_1
XFILLER_6_481 VPWR VGND sg13g2_fill_2
Xhold927 i_snitch.i_snitch_regfile.mem\[141\] VPWR VGND net959 sg13g2_dlygate4sd3_1
XFILLER_103_508 VPWR VGND sg13g2_fill_1
Xhold949 i_snitch.i_snitch_regfile.mem\[58\] VPWR VGND net981 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[211\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2788
+ net2673 VPWR VGND sg13g2_nand2_1
Xhold938 i_snitch.i_snitch_regfile.mem\[220\] VPWR VGND net970 sg13g2_dlygate4sd3_1
Xfanout2690 data_pdata\[13\]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X
+ net2690 VPWR VGND sg13g2_buf_8
XFILLER_85_948 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1 i_snitch.i_snitch_regfile.mem\[56\]_sg13g2_a21oi_1_A1_Y
+ VPWR i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[120\]_sg13g2_nor2_1_A_Y i_snitch.i_snitch_regfile.mem\[88\]_sg13g2_o21ai_1_A1_Y
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2777
+ net2658 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[32\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[32\] VGND sg13g2_inv_1
XFILLER_53_889 VPWR VGND sg13g2_decap_4
XFILLER_25_569 VPWR VGND sg13g2_fill_2
XFILLER_100_35 VPWR VGND sg13g2_decap_8
XFILLER_80_697 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y
+ VPWR VGND net2498 net2418 i_snitch.i_snitch_regfile.mem\[58\]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[3\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[8\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B
+ i_snitch.inst_addr_o\[18\]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X sg13g2_a221oi_1
XFILLER_20_241 VPWR VGND sg13g2_fill_1
XFILLER_21_775 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y VGND VPWR i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_A1
+ net2303 i_snitch.pc_d\[31\] i_snitch.pc_d\[31\]_sg13g2_a21oi_1_Y_B1 sg13g2_a21oi_1
Xi_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[498\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[455\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[455\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net1008 net2460 net2284 VPWR VGND sg13g2_a22oi_1
XFILLER_106_357 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B_sg13g2_nand4_1_Y
+ net2599 net2556 i_snitch.i_snitch_regfile.mem\[35\]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B
+ VPWR VGND net2602 sg13g2_nand4_1
XFILLER_88_720 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q net3284 VGND VPWR i_snitch.i_snitch_regfile.mem\[350\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[350\] clknet_leaf_93_clk sg13g2_dfrbpq_1
Xcnt_q\[2\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y cnt_q\[2\]_sg13g2_a22oi_1_B2_Y state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1
+ net449 cnt_q\[2\]_sg13g2_dfrbpq_1_Q_D VPWR VGND sg13g2_nor3_1
Xi_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A VPWR i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y
+ i_snitch.i_snitch_regfile.mem\[265\] VGND sg13g2_inv_1
XFILLER_0_646 VPWR VGND sg13g2_decap_8
XFILLER_87_252 VPWR VGND sg13g2_decap_4
XFILLER_76_948 VPWR VGND sg13g2_fill_1
XFILLER_47_127 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[437\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
XFILLER_85_69 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1
+ net88 i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[189\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2774
+ net2653 VPWR VGND sg13g2_nand2_1
Xi_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2
+ data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_Y VPWR i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y
+ VGND i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1
+ sg13g2_o21ai_1
XFILLER_28_396 VPWR VGND sg13g2_fill_2
XFILLER_71_675 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q net3207 VGND VPWR i_snitch.i_snitch_regfile.mem\[179\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[179\] clknet_leaf_121_clk sg13g2_dfrbpq_1
Xi_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[242\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2876
+ net2675 VPWR VGND sg13g2_nand2_1
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_34_51 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y VPWR VGND
+ net2477 i_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1
+ net2441 net2789 i_snitch.i_snitch_regfile.mem\[195\]_sg13g2_dfrbpq_1_Q_D net2909
+ sg13g2_a221oi_1
Xi_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2
+ net2507 i_snitch.sb_d\[8\]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nor4_1_Y
+ net3083 net3077 net3079 i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C
+ VGND VPWR net3081 sg13g2_nor4_2
Xi_snitch.inst_addr_o\[10\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[10\]
+ i_snitch.inst_addr_o\[10\] clknet_leaf_53_clk sg13g2_dfrbpq_2
XFILLER_4_941 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[89\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2
+ VGND net2490 i_snitch.i_snitch_regfile.mem\[40\]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X
+ sg13g2_o21ai_1
Xi_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y i_snitch.sb_d\[15\]_sg13g2_o21ai_1_Y_A2
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_snitch.gpr_waddr\[5\]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y
+ VPWR VGND sg13g2_nand2_2
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2794
+ net2660 VPWR VGND sg13g2_nand2_1
XFILLER_94_701 VPWR VGND sg13g2_decap_8
XFILLER_67_915 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B net2820 i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_X
+ i_snitch.i_snitch_regfile.mem\[143\]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y VPWR VGND
+ sg13g2_nor2_1
XFILLER_39_617 VPWR VGND sg13g2_fill_2
XFILLER_38_105 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A
+ i_snitch.sb_d\[12\]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N
+ VPWR VGND sg13g2_nand2b_1
Xi_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1
+ net2554 i_snitch.pc_d\[28\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2
+ VPWR VGND sg13g2_mux2_1
XFILLER_19_363 VPWR VGND sg13g2_decap_4
XFILLER_35_812 VPWR VGND sg13g2_fill_2
XFILLER_74_491 VPWR VGND sg13g2_decap_8
XFILLER_74_480 VPWR VGND sg13g2_fill_1
XFILLER_90_973 VPWR VGND sg13g2_decap_8
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[32\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2298 net1330 net2495 net1217 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[475\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[475\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2372 net826 net2460 net2252 VPWR VGND sg13g2_a22oi_1
XFILLER_15_580 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y
+ i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B VPWR
+ VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[346\]_sg13g2_a22oi_1_B2_Y
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q net3283 VGND VPWR i_snitch.i_snitch_regfile.mem\[370\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[370\] clknet_leaf_91_clk sg13g2_dfrbpq_1
Xdata_pdata\[18\]_sg13g2_mux2_1_A1 rsp_data_q\[18\] net749 net3049 data_pdata\[18\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q
+ net3196 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[17\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
Xhold702 data_pdata\[1\] VPWR VGND net734 sg13g2_dlygate4sd3_1
Xhold746 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[29\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net778 sg13g2_dlygate4sd3_1
Xhold713 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[19\] VPWR
+ VGND net745 sg13g2_dlygate4sd3_1
Xhold724 i_snitch.i_snitch_regfile.mem\[223\] VPWR VGND net756 sg13g2_dlygate4sd3_1
Xhold735 i_snitch.i_snitch_regfile.mem\[145\] VPWR VGND net767 sg13g2_dlygate4sd3_1
XFILLER_89_539 VPWR VGND sg13g2_decap_8
Xrsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y VPWR rsp_data_q\[14\]_sg13g2_dfrbpq_1_Q_D
+ net1298 VGND sg13g2_inv_1
Xhold779 i_snitch.i_snitch_regfile.mem\[268\] VPWR VGND net811 sg13g2_dlygate4sd3_1
Xhold757 i_snitch.i_snitch_regfile.mem\[479\] VPWR VGND net789 sg13g2_dlygate4sd3_1
Xhold768 i_snitch.i_snitch_regfile.mem\[393\] VPWR VGND net800 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y
+ i_snitch.i_snitch_regfile.mem\[161\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B net2443
+ net2514 net2902 net2773 VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[48\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2768
+ net2667 VPWR VGND sg13g2_nand2_1
Xi_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q net3210 VGND VPWR i_snitch.i_snitch_regfile.mem\[199\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[199\] clknet_leaf_119_clk sg13g2_dfrbpq_1
XFILLER_29_127 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[366\]_sg13g2_o21ai_1_A1 net2970 VPWR i_snitch.i_snitch_regfile.mem\[366\]_sg13g2_o21ai_1_A1_Y
+ VGND i_snitch.i_snitch_regfile.mem\[366\] net2805 sg13g2_o21ai_1
Xi_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y
+ i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B
+ VGND net3077 i_snitch.i_snitch_lsu.metadata_q\[4\]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
Xi_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q net3212 VGND VPWR i_snitch.i_snitch_regfile.mem\[505\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[505\] clknet_leaf_115_clk sg13g2_dfrbpq_1
XFILLER_38_672 VPWR VGND sg13g2_fill_1
XFILLER_72_439 VPWR VGND sg13g2_fill_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_nand2_1_A_Y
+ VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[43\]_sg13g2_dfrbpq_1_Q_D
+ VGND i_req_register.data_o\[43\]_sg13g2_o21ai_1_Y_A2 net2619 sg13g2_o21ai_1
XFILLER_81_984 VPWR VGND sg13g2_decap_8
XFILLER_80_450 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C i_req_arb.data_i\[42\]_sg13g2_inv_1_A_Y
+ net2302 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1 i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C_Y
+ VPWR VGND sg13g2_nor3_1
XFILLER_41_804 VPWR VGND sg13g2_decap_8
XFILLER_41_815 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q net3299 VGND VPWR i_snitch.i_snitch_regfile.mem\[47\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[47\] clknet_leaf_63_clk sg13g2_dfrbpq_2
XFILLER_41_859 VPWR VGND sg13g2_decap_8
Xi_snitch.inst_addr_o\[30\]_sg13g2_dfrbpq_1_Q net3312 VGND VPWR i_snitch.pc_d\[30\]
+ i_snitch.inst_addr_o\[30\] clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_40_347 VPWR VGND sg13g2_fill_1
XFILLER_21_572 VPWR VGND sg13g2_decap_4
Xi_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_A2
+ VGND VPWR i_snitch.i_snitch_regfile.mem\[159\]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B_Y
+ i_snitch.pc_d\[12\]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[64\]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y
+ net2700 sg13g2_a21oi_2
XFILLER_106_154 VPWR VGND sg13g2_decap_8
XFILLER_96_35 VPWR VGND sg13g2_decap_8
XFILLER_0_421 VPWR VGND sg13g2_decap_4
XFILLER_1_944 VPWR VGND sg13g2_decap_8
XFILLER_103_872 VPWR VGND sg13g2_decap_8
XFILLER_0_454 VPWR VGND sg13g2_decap_8
XFILLER_102_371 VPWR VGND sg13g2_decap_8
XFILLER_76_723 VPWR VGND sg13g2_decap_4
XFILLER_49_948 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[495\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[495\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ net2368 net1001 net2678 net2859 VPWR VGND sg13g2_a22oi_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[31\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2
+ i_snitch.i_snitch_regfile.mem\[265\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y
+ net2530 i_snitch.i_snitch_regfile.mem\[65\]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y
+ net2479 VPWR VGND sg13g2_a22oi_1
XFILLER_91_704 VPWR VGND sg13g2_fill_1
XFILLER_91_737 VPWR VGND sg13g2_decap_8
XFILLER_63_428 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q net3291 VGND VPWR i_snitch.i_snitch_regfile.mem\[390\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[390\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_29_672 VPWR VGND sg13g2_fill_2
XFILLER_17_834 VPWR VGND sg13g2_decap_8
Xdata_pdata\[5\]_sg13g2_nor2_1_B net3157 data_pdata\[5\] data_pdata\[5\]_sg13g2_nor2_1_B_Y
+ VPWR VGND sg13g2_nor2_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q
+ net3228 VGND VPWR i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\]_sg13g2_dfrbpq_1_Q_D
+ i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[37\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
XFILLER_44_675 VPWR VGND sg13g2_fill_1
XFILLER_71_472 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1 VGND VPWR
+ i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y net2840 i_snitch.i_snitch_regfile.mem\[325\]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y
+ i_snitch.i_snitch_regfile.mem\[357\]_sg13g2_o21ai_1_A1_Y sg13g2_a21oi_1
XFILLER_32_837 VPWR VGND sg13g2_decap_4
Xi_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A
+ net44 net2718 i_req_arb.gen_arbiter.req_d\[1\]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X
+ VPWR VGND sg13g2_and2_1
XFILLER_77_7 VPWR VGND sg13g2_fill_2
XFILLER_8_554 VPWR VGND sg13g2_decap_4
XFILLER_40_892 VPWR VGND sg13g2_fill_1
XFILLER_99_804 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1
+ VPWR i_snitch.i_snitch_regfile.mem\[459\]_sg13g2_dfrbpq_1_Q_D VGND net2280 net2377
+ sg13g2_o21ai_1
XFILLER_6_77 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[314\]_sg13g2_a22oi_1_A1 i_snitch.i_snitch_regfile.mem\[314\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2430 net2255 net2316 net1205 VPWR VGND sg13g2_a22oi_1
Xstrb_reg_q\[6\]_sg13g2_nand2_1_A strb_reg_q\[6\]_sg13g2_nand2_1_A_Y net442 net3043
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A
+ i_snitch.pc_d\[7\]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_2
XFILLER_66_200 VPWR VGND sg13g2_decap_4
XFILLER_6_1026 VPWR VGND sg13g2_fill_2
XFILLER_94_542 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_mux2_1_A1
+ net998 net665 net68 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[5\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND sg13g2_mux2_1
Xi_snitch.i_snitch_regfile.mem\[67\]_sg13g2_dfrbpq_1_Q net3273 VGND VPWR i_snitch.i_snitch_regfile.mem\[67\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[67\] clknet_leaf_100_clk sg13g2_dfrbpq_1
Xrebuffer27 i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A
+ net59 VPWR VGND sg13g2_buf_1
Xrebuffer16 i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y
+ net48 VPWR VGND sg13g2_buf_2
XFILLER_48_981 VPWR VGND sg13g2_fill_2
Xi_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[461\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2290
+ net2461 VPWR VGND sg13g2_nand2_1
Xrebuffer38 net40 net70 VPWR VGND sg13g2_buf_2
Xrebuffer49 i_snitch.i_snitch_regfile.mem\[129\]_sg13g2_a22oi_1_A1_A2 net81 VPWR VGND
+ sg13g2_buf_8
XFILLER_62_450 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[315\]_sg13g2_a21oi_1_A1 VGND VPWR i_snitch.i_snitch_regfile.mem\[315\]
+ net2999 i_snitch.i_snitch_regfile.mem\[315\]_sg13g2_a21oi_1_A1_Y net2973 sg13g2_a21oi_1
XFILLER_22_314 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[5\]_sg13g2_nor2_1_B_A i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B
+ i_snitch.pc_d\[6\]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A
+ VPWR i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A_Y
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1
+ VGND sg13g2_inv_1
Xi_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2 VPWR
+ VGND i_snitch.i_snitch_regfile.mem\[511\]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y net2957
+ i_snitch.i_snitch_regfile.mem\[415\]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y net2969
+ i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y i_snitch.i_snitch_regfile.mem\[287\]_sg13g2_mux4_1_A0_1_X
+ sg13g2_a221oi_1
Xdata_pdata\[9\]_sg13g2_nand2b_1_B data_pdata\[9\]_sg13g2_nand2b_1_B_Y data_pdata\[9\]
+ net3157 VPWR VGND sg13g2_nand2b_1
Xhold510 shift_reg_q\[22\]_sg13g2_dfrbpq_1_Q_D VPWR VGND net542 sg13g2_dlygate4sd3_1
Xhold521 i_snitch.wake_up_q\[1\] VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold554 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[7\] VPWR
+ VGND net586 sg13g2_dlygate4sd3_1
Xhold532 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\] VPWR
+ VGND net564 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2
+ i_snitch.pc_d\[17\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A net41
+ VPWR VGND sg13g2_xnor2_1
XFILLER_2_719 VPWR VGND sg13g2_decap_8
Xhold543 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[15\]_sg13g2_dfrbpq_1_Q_D
+ VPWR VGND net575 sg13g2_dlygate4sd3_1
XFILLER_104_625 VPWR VGND sg13g2_fill_2
XFILLER_89_336 VPWR VGND sg13g2_fill_1
Xhold576 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[30\] VPWR
+ VGND net608 sg13g2_dlygate4sd3_1
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C net2312 i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1
+ i_snitch.pc_d\[2\]_sg13g2_nor2_1_B_A i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y
+ VPWR VGND sg13g2_nand3_1
Xhold565 i_snitch.i_snitch_regfile.mem\[415\] VPWR VGND net597 sg13g2_dlygate4sd3_1
Xhold587 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[3\] VPWR
+ VGND net619 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[103\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xhold598 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[13\] VPWR
+ VGND net630 sg13g2_dlygate4sd3_1
XFILLER_106_56 VPWR VGND sg13g2_decap_8
XFILLER_103_168 VPWR VGND sg13g2_decap_8
XFILLER_98_892 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[13\]_sg13g2_a21o_1_X net2305 net1375 i_snitch.pc_d\[13\]_sg13g2_a21o_1_X_B1
+ i_snitch.pc_d\[13\] VPWR VGND sg13g2_a21o_1
XFILLER_58_734 VPWR VGND sg13g2_decap_8
XFILLER_58_712 VPWR VGND sg13g2_fill_1
Xhold1232 rsp_data_q\[4\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A VPWR VGND net1264 sg13g2_dlygate4sd3_1
Xhold1210 i_snitch.inst_addr_o\[21\] VPWR VGND net1242 sg13g2_dlygate4sd3_1
Xhold1221 i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[40\] VPWR
+ VGND net1253 sg13g2_dlygate4sd3_1
Xhold1243 i_snitch.i_snitch_regfile.mem\[176\] VPWR VGND net1275 sg13g2_dlygate4sd3_1
Xi_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[391\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y
+ net123 i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0
+ i_snitch.pc_d\[5\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1
+ VPWR VGND sg13g2_nor2_1
XFILLER_100_875 VPWR VGND sg13g2_decap_8
Xhold1265 rsp_data_q\[14\] VPWR VGND net1297 sg13g2_dlygate4sd3_1
XFILLER_57_277 VPWR VGND sg13g2_fill_2
Xhold1276 i_snitch.i_snitch_regfile.mem\[413\] VPWR VGND net1308 sg13g2_dlygate4sd3_1
Xhold1254 i_snitch.i_snitch_regfile.mem\[130\] VPWR VGND net1286 sg13g2_dlygate4sd3_1
Xhold1287 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q VPWR VGND
+ net1319 sg13g2_dlygate4sd3_1
Xhold1298 rsp_data_q\[26\] VPWR VGND net1330 sg13g2_dlygate4sd3_1
Xi_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]_sg13g2_nand2_1_B
+ i_req_register.data_o\[45\]_sg13g2_o21ai_1_Y_B1 net3169 i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[45\]
+ VPWR VGND sg13g2_nand2_1
Xdata_pdata\[8\]_sg13g2_dfrbpq_1_Q net3228 VGND VPWR net1148 data_pdata\[8\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
XFILLER_17_119 VPWR VGND sg13g2_fill_1
XFILLER_72_247 VPWR VGND sg13g2_fill_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A
+ net2933 net2919 i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[19\]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y
+ VPWR VGND sg13g2_nand3_1
Xrsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y rsp_data_q\[20\]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A
+ net3058 net907 net3063 rsp_data_q\[16\] VPWR VGND sg13g2_a22oi_1
Xi_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A i_snitch.i_snitch_regfile.mem\[330\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ VPWR VGND sg13g2_nand2_1
Xi_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y
+ VPWR VGND net2548 i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D
+ i_snitch.i_snitch_regfile.mem\[407\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C
+ i_snitch.pc_d\[23\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2
+ sg13g2_a221oi_1
XFILLER_40_199 VPWR VGND sg13g2_decap_8
Xi_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y
+ i_snitch.pc_d\[2\]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B
+ VPWR VGND sg13g2_xnor2_1
Xi_snitch.i_snitch_regfile.mem\[334\]_sg13g2_a22oi_1_B2 i_snitch.i_snitch_regfile.mem\[334\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B
+ net2405 net947 net2687 net2798 VPWR VGND sg13g2_a22oi_1
XFILLER_103_0 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q net3323 VGND VPWR i_snitch.i_snitch_regfile.mem\[87\]_sg13g2_dfrbpq_1_Q_D
+ i_snitch.i_snitch_regfile.mem\[87\] clknet_leaf_60_clk sg13g2_dfrbpq_1
XFILLER_1_741 VPWR VGND sg13g2_decap_8
XFILLER_89_881 VPWR VGND sg13g2_decap_8
XFILLER_49_745 VPWR VGND sg13g2_fill_1
XFILLER_48_222 VPWR VGND sg13g2_fill_1
Xi_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y
+ net2543 VPWR i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1
+ VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y
+ i_snitch.pc_d\[10\]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2
+ sg13g2_o21ai_1
XFILLER_91_534 VPWR VGND sg13g2_fill_2
XFILLER_64_748 VPWR VGND sg13g2_fill_1
XFILLER_91_556 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A_sg13g2_nor2_1_Y
+ i_snitch.pc_d\[9\]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A
+ net2599 i_snitch.pc_d\[18\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A
+ VPWR VGND sg13g2_nor2_1
Xi_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_inv_1_A
+ i_snitch.pc_d\[29\]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A
+ i_snitch.i_snitch_regfile.mem\[445\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ VPWR VGND sg13g2_inv_2
XFILLER_60_943 VPWR VGND sg13g2_decap_4
XFILLER_44_494 VPWR VGND sg13g2_fill_1
Xi_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y
+ i_snitch.i_snitch_regfile.mem\[90\]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A net2782
+ net2660 VPWR VGND sg13g2_nand2_1
XFILLER_31_133 VPWR VGND sg13g2_decap_8
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1
+ VPWR VGND i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[2\]_sg13g2_nand2_1_B_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[0\]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[1\]_sg13g2_nand3b_1_B_Y
+ sg13g2_a221oi_1
Xi_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1
+ i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N_Y
+ VPWR i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q\[21\]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y
+ VGND net3183 i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q\[21\]
+ sg13g2_o21ai_1
XFILLER_31_144 VPWR VGND sg13g2_fill_2
XFILLER_31_177 VPWR VGND sg13g2_fill_2
Xi_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_D
+ i_snitch.pc_d\[8\]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C_Y i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_C
+ i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y VGND VPWR i_snitch.pc_d\[11\]_sg13g2_a21o_1_A2_X
+ sg13g2_nor4_2
XFILLER_9_841 VPWR VGND sg13g2_fill_1
XFILLER_100_105 VPWR VGND sg13g2_decap_8
Xi_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X
+ i_snitch.i_snitch_regfile.mem\[261\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C
+ i_snitch.i_snitch_regfile.mem\[394\]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y
+ i_snitch.i_snitch_regfile.mem\[427\]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2
+ VPWR VGND sg13g2_nand3_1
.ends

