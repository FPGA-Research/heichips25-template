module heichips25_snitch_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \cnt_q[0] ;
 wire \cnt_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \cnt_q[1] ;
 wire \cnt_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \cnt_q[2] ;
 wire \cnt_q[2]_sg13g2_a21oi_1_B1_Y ;
 wire \cnt_q[2]_sg13g2_a22oi_1_B2_A2 ;
 wire \cnt_q[2]_sg13g2_a22oi_1_B2_B1 ;
 wire \cnt_q[2]_sg13g2_a22oi_1_B2_Y ;
 wire \cnt_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \cnt_q[2]_sg13g2_nand3_1_A_Y ;
 wire \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X ;
 wire \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ;
 wire \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[0] ;
 wire \data_pdata[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[0]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[0]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[10] ;
 wire \data_pdata[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[10]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ;
 wire \data_pdata[10]_sg13g2_nor2b_1_A_Y ;
 wire \data_pdata[11] ;
 wire \data_pdata[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[11]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ;
 wire \data_pdata[11]_sg13g2_nor2b_1_A_Y ;
 wire \data_pdata[12] ;
 wire \data_pdata[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[12]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ;
 wire \data_pdata[12]_sg13g2_nor2b_1_A_Y ;
 wire \data_pdata[13] ;
 wire \data_pdata[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[13]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ;
 wire \data_pdata[13]_sg13g2_nor2b_1_A_Y ;
 wire \data_pdata[14] ;
 wire \data_pdata[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[14]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ;
 wire \data_pdata[15] ;
 wire \data_pdata[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[15]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y ;
 wire \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ;
 wire \data_pdata[16] ;
 wire \data_pdata[16]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[16]_sg13g2_nor2b_1_B_N_Y ;
 wire \data_pdata[17] ;
 wire \data_pdata[17]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[17]_sg13g2_nor2b_1_B_N_Y ;
 wire \data_pdata[18] ;
 wire \data_pdata[18]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[18]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ;
 wire \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ;
 wire \data_pdata[19] ;
 wire \data_pdata[19]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[19]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ;
 wire \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ;
 wire \data_pdata[1] ;
 wire \data_pdata[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[1]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[1]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[20] ;
 wire \data_pdata[20]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[20]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ;
 wire \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ;
 wire \data_pdata[21] ;
 wire \data_pdata[21]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[21]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y ;
 wire \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[22] ;
 wire \data_pdata[22]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[22]_sg13g2_nor2b_1_B_N_Y ;
 wire \data_pdata[23] ;
 wire \data_pdata[23]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[23]_sg13g2_nor2b_1_B_N_Y ;
 wire \data_pdata[24] ;
 wire \data_pdata[24]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[24]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[24]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[25] ;
 wire \data_pdata[25]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[25]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[25]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[26] ;
 wire \data_pdata[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[26]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[26]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[27] ;
 wire \data_pdata[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[27]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[27]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[28] ;
 wire \data_pdata[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[28]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[28]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[29] ;
 wire \data_pdata[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[29]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[29]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[2] ;
 wire \data_pdata[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[2]_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[2]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ;
 wire \data_pdata[30] ;
 wire \data_pdata[30]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[30]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[30]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[31] ;
 wire \data_pdata[31]_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[31]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[31]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ;
 wire \data_pdata[3] ;
 wire \data_pdata[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[3]_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[3]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ;
 wire \data_pdata[4] ;
 wire \data_pdata[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[4]_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[4]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ;
 wire \data_pdata[5] ;
 wire \data_pdata[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[5]_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ;
 wire \data_pdata[6] ;
 wire \data_pdata[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[6]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[6]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[7] ;
 wire \data_pdata[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[7]_sg13g2_mux2_1_A0_X ;
 wire \data_pdata[7]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \data_pdata[8] ;
 wire \data_pdata[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[8]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ;
 wire \data_pdata[9] ;
 wire \data_pdata[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \data_pdata[9]_sg13g2_nand2b_1_B_Y ;
 wire \data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ;
 wire \data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ;
 wire data_pvalid;
 wire data_pvalid_sg13g2_dfrbpq_1_Q_D;
 wire data_pvalid_sg13g2_nand2b_1_B_Y;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_X;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D;
 wire data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y;
 wire data_pvalid_sg13g2_nor2_1_A_B;
 wire data_pvalid_sg13g2_nor2_1_A_Y;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_B1;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D_X;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A_Y;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B;
 wire data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y;
 wire data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A ;
 wire \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B ;
 wire \i_req_arb.data_i[37] ;
 wire \i_req_arb.data_i[38] ;
 wire \i_req_arb.data_i[39] ;
 wire \i_req_arb.data_i[40] ;
 wire \i_req_arb.data_i[41] ;
 wire \i_req_arb.data_i[42] ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2 ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1 ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ;
 wire \i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ;
 wire \i_req_arb.data_i[43] ;
 wire \i_req_arb.data_i[44] ;
 wire \i_req_arb.data_i[44]_sg13g2_a21o_1_B1_X ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1 ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A_Y ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[0] ;
 wire \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[1] ;
 wire \i_req_arb.gen_arbiter.req_d[1] ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_o21ai_1_A2_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_A ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_C ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1 ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X ;
 wire \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y ;
 wire \i_req_arb.gen_arbiter.rr_q ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2 ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1 ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B_X ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y ;
 wire \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A_X ;
 wire \i_req_register.data_o[38] ;
 wire \i_req_register.data_o[39] ;
 wire \i_req_register.data_o[39]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.data_o[39]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.data_o[40] ;
 wire \i_req_register.data_o[41] ;
 wire \i_req_register.data_o[41]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.data_o[41]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.data_o[42] ;
 wire \i_req_register.data_o[43] ;
 wire \i_req_register.data_o[43]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.data_o[43]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.data_o[44] ;
 wire \i_req_register.data_o[44]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.data_o[44]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.data_o[45] ;
 wire \i_req_register.data_o[45]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.data_o[45]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.data_o[5] ;
 wire \i_req_register.data_o[5]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_nand2_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_nand2_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_nand2_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_nand2_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1_1_X ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q ;
 wire \i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.consec_pc[0] ;
 wire \i_snitch.consec_pc[0]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.gpr_waddr[4] ;
 wire \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.gpr_waddr[5] ;
 wire \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ;
 wire \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.gpr_waddr[6] ;
 wire \i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.gpr_waddr[7] ;
 wire \i_snitch.gpr_waddr[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_d ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_q ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_or2_1_A_X ;
 wire \i_snitch.i_snitch_lsu.metadata_q[1] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[2] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[3] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_lsu.metadata_q[9] ;
 wire \i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[100] ;
 wire \i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[100]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[101] ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[102] ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[102]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[103] ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[103]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[104] ;
 wire \i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[104]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[105] ;
 wire \i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[106] ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[107] ;
 wire \i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[108] ;
 wire \i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[109] ;
 wire \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[110] ;
 wire \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[111] ;
 wire \i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[111]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[112] ;
 wire \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[113] ;
 wire \i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[114] ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[115] ;
 wire \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[116] ;
 wire \i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[117] ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[118] ;
 wire \i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[119] ;
 wire \i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[120] ;
 wire \i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[121] ;
 wire \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[122] ;
 wire \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[123] ;
 wire \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[124] ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[125] ;
 wire \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[126] ;
 wire \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[127] ;
 wire \i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[128] ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[129] ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[130] ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[131] ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[132] ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[133] ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[134] ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[135] ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[136] ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[137] ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[138] ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[139] ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[140] ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[141] ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[142] ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[143] ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[144] ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[145] ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[146] ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[147] ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[148] ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[149] ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[150] ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2 ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[151] ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[152] ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[153] ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[154] ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[155] ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[156] ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[157] ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[158] ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[159] ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[160] ;
 wire \i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[161] ;
 wire \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[161]_sg13g2_nand2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[162] ;
 wire \i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[163] ;
 wire \i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[164] ;
 wire \i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[165] ;
 wire \i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[166] ;
 wire \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[167] ;
 wire \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[168] ;
 wire \i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[169] ;
 wire \i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[170] ;
 wire \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[171] ;
 wire \i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[172] ;
 wire \i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[173] ;
 wire \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[174] ;
 wire \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[175] ;
 wire \i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[176] ;
 wire \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[177] ;
 wire \i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[178] ;
 wire \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[179] ;
 wire \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[180] ;
 wire \i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[181] ;
 wire \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[182] ;
 wire \i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[183] ;
 wire \i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[184] ;
 wire \i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[185] ;
 wire \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[186] ;
 wire \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[187] ;
 wire \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[188] ;
 wire \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[189] ;
 wire \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[190] ;
 wire \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[191] ;
 wire \i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[192] ;
 wire \i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[193] ;
 wire \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[194] ;
 wire \i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[195] ;
 wire \i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[196] ;
 wire \i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[197] ;
 wire \i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[198] ;
 wire \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[199] ;
 wire \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[200] ;
 wire \i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[201] ;
 wire \i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[202] ;
 wire \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[203] ;
 wire \i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[204] ;
 wire \i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[205] ;
 wire \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[206] ;
 wire \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[207] ;
 wire \i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[208] ;
 wire \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[209] ;
 wire \i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[210] ;
 wire \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[211] ;
 wire \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[212] ;
 wire \i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[213] ;
 wire \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[214] ;
 wire \i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[215] ;
 wire \i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[216] ;
 wire \i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[217] ;
 wire \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[218] ;
 wire \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[219] ;
 wire \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[220] ;
 wire \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[221] ;
 wire \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[222] ;
 wire \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[223] ;
 wire \i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[224] ;
 wire \i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[225] ;
 wire \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[226] ;
 wire \i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[227] ;
 wire \i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[228] ;
 wire \i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[229] ;
 wire \i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[230] ;
 wire \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[231] ;
 wire \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[232] ;
 wire \i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[233] ;
 wire \i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[234] ;
 wire \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[235] ;
 wire \i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[236] ;
 wire \i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[237] ;
 wire \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[238] ;
 wire \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[239] ;
 wire \i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[240] ;
 wire \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[241] ;
 wire \i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[242] ;
 wire \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[243] ;
 wire \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[244] ;
 wire \i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[245] ;
 wire \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[246] ;
 wire \i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[247] ;
 wire \i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[248] ;
 wire \i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[249] ;
 wire \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[250] ;
 wire \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[251] ;
 wire \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[252] ;
 wire \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[253] ;
 wire \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[254] ;
 wire \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[255] ;
 wire \i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[256] ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[257] ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[258] ;
 wire \i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[259] ;
 wire \i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[260] ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[261] ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X ;
 wire \i_snitch.i_snitch_regfile.mem[262] ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[263] ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[263]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[264] ;
 wire \i_snitch.i_snitch_regfile.mem[264]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[264]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265] ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[266] ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[267] ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[268] ;
 wire \i_snitch.i_snitch_regfile.mem[268]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[268]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269] ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270] ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[271] ;
 wire \i_snitch.i_snitch_regfile.mem[271]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[271]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[272] ;
 wire \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[272]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[272]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273] ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[274] ;
 wire \i_snitch.i_snitch_regfile.mem[274]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[274]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[275] ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[276] ;
 wire \i_snitch.i_snitch_regfile.mem[276]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[276]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[277] ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[278] ;
 wire \i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[278]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[279] ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[280] ;
 wire \i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[280]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[280]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281] ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[282] ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283] ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[284] ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[284]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[285] ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[285]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286] ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[287] ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[288] ;
 wire \i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[288]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[289] ;
 wire \i_snitch.i_snitch_regfile.mem[289]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[290] ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[291] ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B ;
 wire \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[292] ;
 wire \i_snitch.i_snitch_regfile.mem[292]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[293] ;
 wire \i_snitch.i_snitch_regfile.mem[293]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[294] ;
 wire \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[294]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[295] ;
 wire \i_snitch.i_snitch_regfile.mem[295]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[296] ;
 wire \i_snitch.i_snitch_regfile.mem[296]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[296]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[297] ;
 wire \i_snitch.i_snitch_regfile.mem[297]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[297]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[298] ;
 wire \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[298]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[299] ;
 wire \i_snitch.i_snitch_regfile.mem[299]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[300] ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[300]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[301] ;
 wire \i_snitch.i_snitch_regfile.mem[301]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[301]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[302] ;
 wire \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[302]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[302]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[303] ;
 wire \i_snitch.i_snitch_regfile.mem[303]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[303]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304] ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[305] ;
 wire \i_snitch.i_snitch_regfile.mem[305]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[305]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[306] ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[306]_sg13g2_nand2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[307] ;
 wire \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[307]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308] ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[308]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[309] ;
 wire \i_snitch.i_snitch_regfile.mem[309]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[309]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[310] ;
 wire \i_snitch.i_snitch_regfile.mem[310]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[311] ;
 wire \i_snitch.i_snitch_regfile.mem[311]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[312] ;
 wire \i_snitch.i_snitch_regfile.mem[312]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[313] ;
 wire \i_snitch.i_snitch_regfile.mem[313]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[313]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[314] ;
 wire \i_snitch.i_snitch_regfile.mem[314]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[314]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[315] ;
 wire \i_snitch.i_snitch_regfile.mem[315]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[315]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[316] ;
 wire \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[317] ;
 wire \i_snitch.i_snitch_regfile.mem[317]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[318] ;
 wire \i_snitch.i_snitch_regfile.mem[318]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[318]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[319] ;
 wire \i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[320] ;
 wire \i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[320]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[321] ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[321]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[322] ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[323] ;
 wire \i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[323]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[324] ;
 wire \i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[325] ;
 wire \i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[326] ;
 wire \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[326]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[327] ;
 wire \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[328] ;
 wire \i_snitch.i_snitch_regfile.mem[328]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[328]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[329] ;
 wire \i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[329]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32] ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[330] ;
 wire \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[330]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[331] ;
 wire \i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[332] ;
 wire \i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[332]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[333] ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[333]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[334] ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[334]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[335] ;
 wire \i_snitch.i_snitch_regfile.mem[335]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[335]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[336] ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[336]_sg13g2_nand2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[337] ;
 wire \i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[337]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[338] ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[339] ;
 wire \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[339]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[33] ;
 wire \i_snitch.i_snitch_regfile.mem[33]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[33]_sg13g2_nand2_1_A_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[340] ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[340]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[341] ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[342] ;
 wire \i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[343] ;
 wire \i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[344] ;
 wire \i_snitch.i_snitch_regfile.mem[344]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[344]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[345] ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[345]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[346] ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[347] ;
 wire \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[347]_sg13g2_nor2b_1_B_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[347]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[348] ;
 wire \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[348]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[349] ;
 wire \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34] ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A_C ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_X ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[34]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[350] ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[350]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[351] ;
 wire \i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[352] ;
 wire \i_snitch.i_snitch_regfile.mem[352]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[353] ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[354] ;
 wire \i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[354]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[354]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[355] ;
 wire \i_snitch.i_snitch_regfile.mem[355]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[356] ;
 wire \i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[356]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[357] ;
 wire \i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[357]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[358] ;
 wire \i_snitch.i_snitch_regfile.mem[358]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[359] ;
 wire \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[359]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35] ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[35]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[360] ;
 wire \i_snitch.i_snitch_regfile.mem[360]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[360]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[361] ;
 wire \i_snitch.i_snitch_regfile.mem[361]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[361]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[362] ;
 wire \i_snitch.i_snitch_regfile.mem[362]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[363] ;
 wire \i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[363]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[364] ;
 wire \i_snitch.i_snitch_regfile.mem[364]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[364]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[365] ;
 wire \i_snitch.i_snitch_regfile.mem[365]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[365]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[366] ;
 wire \i_snitch.i_snitch_regfile.mem[366]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[366]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[367] ;
 wire \i_snitch.i_snitch_regfile.mem[367]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[367]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[368] ;
 wire \i_snitch.i_snitch_regfile.mem[368]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[368]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[369] ;
 wire \i_snitch.i_snitch_regfile.mem[369]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[369]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[36] ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[36]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[370] ;
 wire \i_snitch.i_snitch_regfile.mem[370]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[370]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[371] ;
 wire \i_snitch.i_snitch_regfile.mem[371]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[372] ;
 wire \i_snitch.i_snitch_regfile.mem[372]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[372]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[373] ;
 wire \i_snitch.i_snitch_regfile.mem[373]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[373]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[374] ;
 wire \i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[374]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[375] ;
 wire \i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[375]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[376] ;
 wire \i_snitch.i_snitch_regfile.mem[376]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[376]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[377] ;
 wire \i_snitch.i_snitch_regfile.mem[377]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[377]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[378] ;
 wire \i_snitch.i_snitch_regfile.mem[378]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[378]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[379] ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[37] ;
 wire \i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[37]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[37]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[380] ;
 wire \i_snitch.i_snitch_regfile.mem[380]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[381] ;
 wire \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[381]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[382] ;
 wire \i_snitch.i_snitch_regfile.mem[382]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[382]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[383] ;
 wire \i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[384] ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[385] ;
 wire \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[386] ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[387] ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388] ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[389] ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[38] ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[38]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[390] ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[391] ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[392] ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[393] ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[394] ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[395] ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[395]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[396] ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[397] ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[398] ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[398]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[399] ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[39] ;
 wire \i_snitch.i_snitch_regfile.mem[39]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[39]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[400] ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[401] ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[402] ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[403] ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[403]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[404] ;
 wire \i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[404]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[405] ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[406] ;
 wire \i_snitch.i_snitch_regfile.mem[406]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[406]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407] ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[408] ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[409] ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[40] ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[40]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[410] ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[411] ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[412] ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[413] ;
 wire \i_snitch.i_snitch_regfile.mem[413]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[413]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[414] ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.i_snitch_regfile.mem[415] ;
 wire \i_snitch.i_snitch_regfile.mem[415]_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[415]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[416] ;
 wire \i_snitch.i_snitch_regfile.mem[416]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[417] ;
 wire \i_snitch.i_snitch_regfile.mem[417]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[418] ;
 wire \i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[419] ;
 wire \i_snitch.i_snitch_regfile.mem[419]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[41] ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[420] ;
 wire \i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[421] ;
 wire \i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[421]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[422] ;
 wire \i_snitch.i_snitch_regfile.mem[422]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[423] ;
 wire \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[423]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[424] ;
 wire \i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[425] ;
 wire \i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[426] ;
 wire \i_snitch.i_snitch_regfile.mem[426]_sg13g2_a21o_1_A1_X ;
 wire \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[427] ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ;
 wire \i_snitch.i_snitch_regfile.mem[428] ;
 wire \i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[429] ;
 wire \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[42] ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[430] ;
 wire \i_snitch.i_snitch_regfile.mem[430]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[431] ;
 wire \i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[432] ;
 wire \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[433] ;
 wire \i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[434] ;
 wire \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[435] ;
 wire \i_snitch.i_snitch_regfile.mem[435]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[436] ;
 wire \i_snitch.i_snitch_regfile.mem[436]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[437] ;
 wire \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[438] ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[438]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[439] ;
 wire \i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[439]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[43] ;
 wire \i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[43]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[440] ;
 wire \i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[440]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[441] ;
 wire \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[442] ;
 wire \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[443] ;
 wire \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[444] ;
 wire \i_snitch.i_snitch_regfile.mem[444]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[445] ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[445]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[446] ;
 wire \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[447] ;
 wire \i_snitch.i_snitch_regfile.mem[447]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[447]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[448] ;
 wire \i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[448]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[449] ;
 wire \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[449]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[44] ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[450] ;
 wire \i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[451] ;
 wire \i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[452] ;
 wire \i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[452]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[453] ;
 wire \i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[453]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[454] ;
 wire \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[455] ;
 wire \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[455]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[456] ;
 wire \i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[457] ;
 wire \i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[458] ;
 wire \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[458]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[459] ;
 wire \i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[459]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[45] ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[460] ;
 wire \i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[461] ;
 wire \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[462] ;
 wire \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[463] ;
 wire \i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[464] ;
 wire \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[465] ;
 wire \i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[466] ;
 wire \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[467] ;
 wire \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[468] ;
 wire \i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[469] ;
 wire \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[46] ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[46]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[470] ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[470]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[471] ;
 wire \i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[471]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[472] ;
 wire \i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[473] ;
 wire \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[474] ;
 wire \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[475] ;
 wire \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[476] ;
 wire \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[477] ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[477]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[478] ;
 wire \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[479] ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47] ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[47]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[480] ;
 wire \i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[481] ;
 wire \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[482] ;
 wire \i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[483] ;
 wire \i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[483]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[484] ;
 wire \i_snitch.i_snitch_regfile.mem[484]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[485] ;
 wire \i_snitch.i_snitch_regfile.mem[485]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[486] ;
 wire \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[486]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[487] ;
 wire \i_snitch.i_snitch_regfile.mem[487]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[488] ;
 wire \i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[489] ;
 wire \i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[48] ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[48]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[490] ;
 wire \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[491] ;
 wire \i_snitch.i_snitch_regfile.mem[491]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[492] ;
 wire \i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[493] ;
 wire \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[494] ;
 wire \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[494]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[495] ;
 wire \i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[496] ;
 wire \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[497] ;
 wire \i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[498] ;
 wire \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[499] ;
 wire \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[499]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[49] ;
 wire \i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[49]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[500] ;
 wire \i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[500]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[501] ;
 wire \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[502] ;
 wire \i_snitch.i_snitch_regfile.mem[502]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[502]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[503] ;
 wire \i_snitch.i_snitch_regfile.mem[503]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[504] ;
 wire \i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[504]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[505] ;
 wire \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[506] ;
 wire \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[507] ;
 wire \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[508] ;
 wire \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[508]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[509] ;
 wire \i_snitch.i_snitch_regfile.mem[509]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[509]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[50] ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[510] ;
 wire \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[511] ;
 wire \i_snitch.i_snitch_regfile.mem[511]_sg13g2_a21o_1_A1_X ;
 wire \i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51] ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[52] ;
 wire \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[53] ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[54] ;
 wire \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[55] ;
 wire \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[56] ;
 wire \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[57] ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[57]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[58] ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[58]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[59] ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[60] ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[61] ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[61]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[62] ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63] ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_B ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[64] ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[64]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[65] ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[66] ;
 wire \i_snitch.i_snitch_regfile.mem[66]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[66]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[66]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[66]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[67] ;
 wire \i_snitch.i_snitch_regfile.mem[67]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[67]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[67]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[67]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[68] ;
 wire \i_snitch.i_snitch_regfile.mem[68]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[68]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[68]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[68]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[69] ;
 wire \i_snitch.i_snitch_regfile.mem[69]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[69]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[69]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[69]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[70] ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[71] ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[72] ;
 wire \i_snitch.i_snitch_regfile.mem[72]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[73] ;
 wire \i_snitch.i_snitch_regfile.mem[73]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[73]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[74] ;
 wire \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[74]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[74]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[75] ;
 wire \i_snitch.i_snitch_regfile.mem[75]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[75]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[76] ;
 wire \i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[76]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[76]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[77] ;
 wire \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[77]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[77]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[78] ;
 wire \i_snitch.i_snitch_regfile.mem[78]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[78]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[79] ;
 wire \i_snitch.i_snitch_regfile.mem[79]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[80] ;
 wire \i_snitch.i_snitch_regfile.mem[80]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[80]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[81] ;
 wire \i_snitch.i_snitch_regfile.mem[81]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[81]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[82] ;
 wire \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[82]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[82]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[83] ;
 wire \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[83]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[83]_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[84] ;
 wire \i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[84]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[84]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[85] ;
 wire \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[85]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[85]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[86] ;
 wire \i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[86]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[86]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[87] ;
 wire \i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[87]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[87]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[88] ;
 wire \i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[88]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[88]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[89] ;
 wire \i_snitch.i_snitch_regfile.mem[89]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[89]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[90] ;
 wire \i_snitch.i_snitch_regfile.mem[90]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[90]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[91] ;
 wire \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[91]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[91]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[92] ;
 wire \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[92]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[92]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[93] ;
 wire \i_snitch.i_snitch_regfile.mem[93]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[93]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[94] ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[94]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[95] ;
 wire \i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[95]_sg13g2_mux2_1_A0_X ;
 wire \i_snitch.i_snitch_regfile.mem[95]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[96] ;
 wire \i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[96]_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.i_snitch_regfile.mem[97] ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[98] ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_B ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[99] ;
 wire \i_snitch.i_snitch_regfile.mem[99]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.i_snitch_regfile.mem[99]_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.i_snitch_regfile.mem[99]_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.inst_addr_o[10] ;
 wire \i_snitch.inst_addr_o[11] ;
 wire \i_snitch.inst_addr_o[12] ;
 wire \i_snitch.inst_addr_o[13] ;
 wire \i_snitch.inst_addr_o[14] ;
 wire \i_snitch.inst_addr_o[15] ;
 wire \i_snitch.inst_addr_o[16] ;
 wire \i_snitch.inst_addr_o[17] ;
 wire \i_snitch.inst_addr_o[18] ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1_A1 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N_B ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ;
 wire \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ;
 wire \i_snitch.inst_addr_o[19] ;
 wire \i_snitch.inst_addr_o[1] ;
 wire \i_snitch.inst_addr_o[20] ;
 wire \i_snitch.inst_addr_o[21] ;
 wire \i_snitch.inst_addr_o[22] ;
 wire \i_snitch.inst_addr_o[23] ;
 wire \i_snitch.inst_addr_o[24] ;
 wire \i_snitch.inst_addr_o[25] ;
 wire \i_snitch.inst_addr_o[26] ;
 wire \i_snitch.inst_addr_o[27] ;
 wire \i_snitch.inst_addr_o[28] ;
 wire \i_snitch.inst_addr_o[29] ;
 wire \i_snitch.inst_addr_o[30] ;
 wire \i_snitch.inst_addr_o[31] ;
 wire \i_snitch.pc_d[0] ;
 wire \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[10] ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[11] ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_C ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_D ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B_X ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12] ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_C ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.pc_d[12]_sg13g2_mux2_1_A1_A0 ;
 wire \i_snitch.pc_d[12]_sg13g2_mux2_1_A1_X ;
 wire \i_snitch.pc_d[13] ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_A ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14] ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_C1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B_X ;
 wire \i_snitch.pc_d[15] ;
 wire \i_snitch.pc_d[15]_sg13g2_a21o_1_A2_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X ;
 wire \i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A_X ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[16] ;
 wire \i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_B2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17] ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[18] ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X ;
 wire \i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.pc_d[19] ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[1] ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A_X ;
 wire \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[20] ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[20]_sg13g2_or2_1_B_X ;
 wire \i_snitch.pc_d[20]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[21] ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1_A1 ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[22] ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_inv_1_A_Y ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[22]_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[23] ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_B2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X ;
 wire \i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.pc_d[24] ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X ;
 wire \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C_Y ;
 wire \i_snitch.pc_d[25] ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A_X ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[26] ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[26]_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[27] ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[28] ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[28]_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[29] ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_C ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B_X ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C ;
 wire \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A_Y ;
 wire \i_snitch.pc_d[2] ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ;
 wire \i_snitch.pc_d[2]_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[30] ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[31] ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_A_N ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A_X ;
 wire \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[3] ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[4] ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[5] ;
 wire \i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ;
 wire \i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_B_N ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[6] ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_A ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ;
 wire \i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_B1 ;
 wire \i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[7] ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ;
 wire \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C_Y ;
 wire \i_snitch.pc_d[8] ;
 wire \i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A_X ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_C ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y ;
 wire \i_snitch.pc_d[9] ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1 ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N_Y ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B_X ;
 wire \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[10] ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[11] ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[12] ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[13] ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[14] ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[15] ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[1] ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[2] ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[3] ;
 wire \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ;
 wire \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y ;
 wire \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[4] ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[5] ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[6] ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[7] ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[8] ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[9] ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2 ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1 ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ;
 wire \i_snitch.sb_q[10] ;
 wire \i_snitch.sb_q[11] ;
 wire \i_snitch.sb_q[12] ;
 wire \i_snitch.sb_q[13] ;
 wire \i_snitch.sb_q[14] ;
 wire \i_snitch.sb_q[15] ;
 wire \i_snitch.sb_q[1] ;
 wire \i_snitch.sb_q[2] ;
 wire \i_snitch.sb_q[3] ;
 wire \i_snitch.sb_q[4] ;
 wire \i_snitch.sb_q[5] ;
 wire \i_snitch.sb_q[6] ;
 wire \i_snitch.sb_q[7] ;
 wire \i_snitch.sb_q[8] ;
 wire \i_snitch.sb_q[9] ;
 wire \i_snitch.wake_up_q[0] ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0 ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1 ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B ;
 wire \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.wake_up_q[1] ;
 wire \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2 ;
 wire \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B ;
 wire \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1 ;
 wire \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2 ;
 wire \i_snitch.wake_up_q[2] ;
 wire \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ;
 wire \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ;
 wire \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ;
 wire \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ;
 wire \i_snitch.wake_up_q[2]_sg13g2_nor4_1_D_Y ;
 wire req_data_valid;
 wire req_data_valid_sg13g2_o21ai_1_Y_B1;
 wire \rsp_data_q[0] ;
 wire \rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[10] ;
 wire \rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[11] ;
 wire \rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[12] ;
 wire \rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[13] ;
 wire \rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[14] ;
 wire \rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[15] ;
 wire \rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[16] ;
 wire \rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[17] ;
 wire \rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[18] ;
 wire \rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[19] ;
 wire \rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[1] ;
 wire \rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[20] ;
 wire \rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[21] ;
 wire \rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[22] ;
 wire \rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[23] ;
 wire \rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[24] ;
 wire \rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[25] ;
 wire \rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[26] ;
 wire \rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[27] ;
 wire \rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[28] ;
 wire \rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[29] ;
 wire \rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[2] ;
 wire \rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[30] ;
 wire \rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[31] ;
 wire \rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[3] ;
 wire \rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[4] ;
 wire \rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[5] ;
 wire \rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[6] ;
 wire \rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[7] ;
 wire \rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[8] ;
 wire \rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire \rsp_data_q[9] ;
 wire \rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ;
 wire rsp_data_ready;
 wire rsp_state_d;
 wire rsp_state_q;
 wire rsp_state_q_sg13g2_nor2_1_A_Y;
 wire \shift_reg_q[0] ;
 wire \shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ;
 wire \shift_reg_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[0]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[10] ;
 wire \shift_reg_q[10]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[10]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[10]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[11] ;
 wire \shift_reg_q[11]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[11]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[11]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[12] ;
 wire \shift_reg_q[12]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[12]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[12]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[13] ;
 wire \shift_reg_q[13]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[13]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[13]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[14] ;
 wire \shift_reg_q[14]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[14]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[14]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[15] ;
 wire \shift_reg_q[15]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[15]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[15]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[16] ;
 wire \shift_reg_q[16]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[16]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[16]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[17] ;
 wire \shift_reg_q[17]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[17]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[17]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[18] ;
 wire \shift_reg_q[18]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[18]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[18]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[19] ;
 wire \shift_reg_q[19]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[19]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[19]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[1] ;
 wire \shift_reg_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[1]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[20] ;
 wire \shift_reg_q[20]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[20]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[20]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[21] ;
 wire \shift_reg_q[21]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[21]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[21]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[22] ;
 wire \shift_reg_q[22]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[22]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[22]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[23] ;
 wire \shift_reg_q[23]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[23]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[23]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[24] ;
 wire \shift_reg_q[24]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ;
 wire \shift_reg_q[24]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[25] ;
 wire \shift_reg_q[25]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ;
 wire \shift_reg_q[25]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[26] ;
 wire \shift_reg_q[26]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ;
 wire \shift_reg_q[26]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[27] ;
 wire \shift_reg_q[27]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ;
 wire \shift_reg_q[27]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[2] ;
 wire \shift_reg_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[2]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[3] ;
 wire \shift_reg_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[3]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[4] ;
 wire \shift_reg_q[4]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[4]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[5] ;
 wire \shift_reg_q[5]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[5]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[6] ;
 wire \shift_reg_q[6]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[6]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[7] ;
 wire \shift_reg_q[7]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[7]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[7]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[8] ;
 wire \shift_reg_q[8]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[8]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[8]_sg13g2_nor2_1_A_Y ;
 wire \shift_reg_q[9] ;
 wire \shift_reg_q[9]_sg13g2_a22oi_1_A1_Y ;
 wire \shift_reg_q[9]_sg13g2_dfrbpq_1_Q_D ;
 wire \shift_reg_q[9]_sg13g2_nor2_1_A_Y ;
 wire state;
 wire state_sg13g2_dfrbpq_1_Q_D;
 wire state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1;
 wire state_sg13g2_inv_1_A_Y;
 wire strb_out;
 wire strb_out_sg13g2_inv_1_Y_A;
 wire \strb_reg_q[0] ;
 wire \strb_reg_q[0]_sg13g2_a22oi_1_A1_B1 ;
 wire \strb_reg_q[0]_sg13g2_a22oi_1_A1_B2 ;
 wire \strb_reg_q[0]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[0]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[1] ;
 wire \strb_reg_q[1]_sg13g2_a21oi_1_A1_Y ;
 wire \strb_reg_q[1]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[1]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[2] ;
 wire \strb_reg_q[2]_sg13g2_a21oi_1_A1_B1 ;
 wire \strb_reg_q[2]_sg13g2_a21oi_1_A1_Y ;
 wire \strb_reg_q[2]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[2]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[3] ;
 wire \strb_reg_q[3]_sg13g2_a21oi_1_A1_Y ;
 wire \strb_reg_q[3]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[3]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[4] ;
 wire \strb_reg_q[4]_sg13g2_a21oi_1_A1_B1 ;
 wire \strb_reg_q[4]_sg13g2_a21oi_1_A1_Y ;
 wire \strb_reg_q[4]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[4]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[5] ;
 wire \strb_reg_q[5]_sg13g2_a21oi_1_A1_Y ;
 wire \strb_reg_q[5]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[5]_sg13g2_nor2_1_A_Y ;
 wire \strb_reg_q[6] ;
 wire \strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D ;
 wire \strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ;
 wire \strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ;
 wire \strb_reg_q[6]_sg13g2_nand2_1_A_Y ;
 wire \strb_reg_q[6]_sg13g2_nor2_1_A_Y ;
 wire target_sel_q;
 wire target_sel_q_sg13g2_dfrbpq_1_Q_D;
 wire target_sel_q_sg13g2_nand2_1_B_Y;
 wire target_sel_q_sg13g2_nand2b_1_A_N_Y;
 wire target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y;
 wire target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B;
 wire target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_Y;
 wire target_sel_q_sg13g2_nor2_1_A_B;
 wire target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B;
 wire target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B_Y;
 wire target_sel_q_sg13g2_nor2_1_A_Y;
 wire clknet_leaf_0_clk;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire uio_out_sg13g2_inv_1_Y_1_A;
 wire uio_out_sg13g2_inv_1_Y_2_A;
 wire uio_out_sg13g2_inv_1_Y_3_A;
 wire uio_out_sg13g2_inv_1_Y_A;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net25;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net230;
 wire net310;
 wire net414;
 wire net419;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;

 sg13g2_dfrbpq_2 \cnt_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\cnt_q[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_o21ai_1 \cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net500),
    .A2(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net1),
    .Y(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A2(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B1 ));
 sg13g2_nand2_1 \cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .A(net500),
    .B(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ));
 sg13g2_dfrbpq_2 \cnt_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\cnt_q[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_o21ai_1 \cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ),
    .A2(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_xnor2_1 \cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A(net543),
    .B(net500));
 sg13g2_nand2_1 \cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\cnt_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .A(net543),
    .B(\cnt_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \cnt_q[2]_sg13g2_a21oi_1_B1  (.A1(\cnt_q[1] ),
    .A2(\cnt_q[0] ),
    .Y(\cnt_q[2]_sg13g2_a21oi_1_B1_Y ),
    .B1(net448));
 sg13g2_a22oi_1 \cnt_q[2]_sg13g2_a22oi_1_B2  (.Y(\cnt_q[2]_sg13g2_a22oi_1_B2_Y ),
    .B1(\cnt_q[2]_sg13g2_a22oi_1_B2_B1 ),
    .B2(net448),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(net1));
 sg13g2_nand2_1 \cnt_q[2]_sg13g2_a22oi_1_B2_B1_sg13g2_nand2_1_Y  (.Y(\cnt_q[2]_sg13g2_a22oi_1_B2_B1 ),
    .A(net1),
    .B(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \cnt_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(net450),
    .Q(\cnt_q[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_nor3_1 \cnt_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y  (.A(\cnt_q[2]_sg13g2_a22oi_1_B2_Y ),
    .B(state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1),
    .C(net449),
    .Y(\cnt_q[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand3_1 \cnt_q[2]_sg13g2_nand3_1_A  (.B(net543),
    .C(net500),
    .A(net448),
    .Y(\cnt_q[2]_sg13g2_nand3_1_A_Y ));
 sg13g2_and2_1 \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B  (.A(state),
    .B(\cnt_q[2]_sg13g2_nand3_1_A_Y ),
    .X(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X ));
 sg13g2_nor2_1 \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B  (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ),
    .B(\cnt_q[2]_sg13g2_nand3_1_A_Y ),
    .Y(state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1));
 sg13g2_nand2_2 \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2_1_Y  (.Y(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ),
    .A(net1),
    .B(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ));
 sg13g2_nand2b_2 \cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B  (.Y(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y ),
    .B(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A ),
    .A_N(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \data_pdata[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net685),
    .Q(\data_pdata[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_mux2_1 \data_pdata[0]_sg13g2_mux2_1_A0  (.A0(\data_pdata[0] ),
    .A1(\data_pdata[8] ),
    .S(net3161),
    .X(\data_pdata[0]_sg13g2_mux2_1_A0_X ));
 sg13g2_nor2_1 \data_pdata[0]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B  (.A(net3153),
    .B(\data_pdata[0]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[0]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_mux2_1 \data_pdata[0]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[0] ),
    .A1(net684),
    .S(net3051),
    .X(\data_pdata[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \data_pdata[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(net825),
    .Q(\data_pdata[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_mux2_1 \data_pdata[10]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[10] ),
    .A1(net824),
    .S(net3048),
    .X(\data_pdata[10]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[10]_sg13g2_nand2b_1_B  (.Y(\data_pdata[10]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[10] ),
    .A_N(net3157));
 sg13g2_a22oi_1 \data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[26]_sg13g2_nand2b_1_B_Y ),
    .B2(net3150),
    .A2(\data_pdata[18]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[10]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21o_2 \data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2  (.A2(\data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070),
    .B1(net2714),
    .X(\data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2b_1 \data_pdata[10]_sg13g2_nor2b_1_A  (.A(\data_pdata[10] ),
    .B_N(net3157),
    .Y(\data_pdata[10]_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \data_pdata[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net996),
    .Q(\data_pdata[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_mux2_1 \data_pdata[11]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[11] ),
    .A1(net995),
    .S(net3049),
    .X(\data_pdata[11]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[11]_sg13g2_nand2b_1_B  (.Y(\data_pdata[11]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[11] ),
    .A_N(net3158));
 sg13g2_a22oi_1 \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[27]_sg13g2_nand2b_1_B_Y ),
    .B2(net3151),
    .A2(\data_pdata[19]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[11]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21oi_2 \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.B1(net2714),
    .Y(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070));
 sg13g2_inv_1 \data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A  (.Y(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .A(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ));
 sg13g2_nor2b_1 \data_pdata[11]_sg13g2_nor2b_1_A  (.A(\data_pdata[11] ),
    .B_N(net3158),
    .Y(\data_pdata[11]_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \data_pdata[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net902),
    .Q(\data_pdata[12] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[12]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[12] ),
    .A1(net901),
    .S(net3051),
    .X(\data_pdata[12]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[12]_sg13g2_nand2b_1_B  (.Y(\data_pdata[12]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[12] ),
    .A_N(net3159));
 sg13g2_a22oi_1 \data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[28]_sg13g2_nand2b_1_B_Y ),
    .B2(net3152),
    .A2(\data_pdata[20]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[12]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21o_2 \data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2  (.A2(\data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070),
    .B1(net2714),
    .X(\data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2b_1 \data_pdata[12]_sg13g2_nor2b_1_A  (.A(\data_pdata[12] ),
    .B_N(net3161),
    .Y(\data_pdata[12]_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \data_pdata[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3202),
    .D(net726),
    .Q(\data_pdata[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[13]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[13] ),
    .A1(net725),
    .S(net3049),
    .X(\data_pdata[13]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[13]_sg13g2_nand2b_1_B  (.Y(\data_pdata[13]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[13] ),
    .A_N(net3155));
 sg13g2_a22oi_1 \data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[29]_sg13g2_nand2b_1_B_Y ),
    .B2(net3150),
    .A2(\data_pdata[21]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[13]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21o_2 \data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2  (.A2(\data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070),
    .B1(net2714),
    .X(\data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2b_1 \data_pdata[13]_sg13g2_nor2b_1_A  (.A(\data_pdata[13] ),
    .B_N(net3155),
    .Y(\data_pdata[13]_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \data_pdata[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(net1036),
    .Q(\data_pdata[14] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[14]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[14] ),
    .A1(net1035),
    .S(net3050),
    .X(\data_pdata[14]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[14]_sg13g2_nand2b_1_B  (.Y(\data_pdata[14]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[14] ),
    .A_N(net3162));
 sg13g2_a22oi_1 \data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[30]_sg13g2_nand2b_1_B_Y ),
    .B2(net3154),
    .A2(\data_pdata[22]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[14]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21o_2 \data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2  (.A2(\data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070),
    .B1(net2714),
    .X(\data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_dfrbpq_1 \data_pdata[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net967),
    .Q(\data_pdata[15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[15]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[15] ),
    .A1(net966),
    .S(net3052),
    .X(\data_pdata[15]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[15]_sg13g2_nand2b_1_B  (.Y(\data_pdata[15]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[15] ),
    .A_N(net3160));
 sg13g2_a22oi_1 \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1  (.Y(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y ),
    .B1(\data_pdata[15]_sg13g2_nand2b_1_B_Y ),
    .B2(\data_pdata[23]_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[31]_sg13g2_nand2b_1_B_Y ),
    .A1(net3152));
 sg13g2_a21oi_2 \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2  (.B1(net2714),
    .Y(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y ),
    .A1(net3070));
 sg13g2_inv_2 \data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A  (.Y(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .A(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a21oi_1 \data_pdata[16]_sg13g2_a21oi_1_A2  (.A1(net3159),
    .A2(\data_pdata[16] ),
    .Y(\data_pdata[16]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3152));
 sg13g2_dfrbpq_1 \data_pdata[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net810),
    .Q(\data_pdata[16] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[16]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[16] ),
    .A1(net809),
    .S(net3050),
    .X(\data_pdata[16]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2b_1 \data_pdata[16]_sg13g2_nor2b_1_B_N  (.A(net3159),
    .B_N(\data_pdata[16] ),
    .Y(\data_pdata[16]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_1 \data_pdata[17]_sg13g2_a21oi_1_A2  (.A1(net3155),
    .A2(\data_pdata[17] ),
    .Y(\data_pdata[17]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3149));
 sg13g2_dfrbpq_1 \data_pdata[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net730),
    .Q(\data_pdata[17] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_mux2_1 \data_pdata[17]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[17] ),
    .A1(net729),
    .S(net3052),
    .X(\data_pdata[17]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2b_1 \data_pdata[17]_sg13g2_nor2b_1_B_N  (.A(net3156),
    .B_N(\data_pdata[17] ),
    .Y(\data_pdata[17]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_1 \data_pdata[18]_sg13g2_a21oi_1_A2  (.A1(net3156),
    .A2(\data_pdata[18] ),
    .Y(\data_pdata[18]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3150));
 sg13g2_dfrbpq_1 \data_pdata[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net750),
    .Q(\data_pdata[18] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[18]_sg13g2_mux2_1_A0  (.A0(\data_pdata[18] ),
    .A1(\data_pdata[26] ),
    .S(net3156),
    .X(\data_pdata[18]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_2 \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2  (.B1(\data_pdata[2]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ),
    .Y(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[18]_sg13g2_mux2_1_A0_X ),
    .A1(net3150));
 sg13g2_nand3b_1 \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C  (.B(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .C(\data_pdata[18]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ),
    .A_N(net3150));
 sg13g2_nand2_2 \data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B  (.Y(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .A(net2681),
    .B(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ));
 sg13g2_mux2_1 \data_pdata[18]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[18] ),
    .A1(net749),
    .S(net3049),
    .X(\data_pdata[18]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \data_pdata[19]_sg13g2_a21oi_1_A2  (.A1(net3158),
    .A2(\data_pdata[19] ),
    .Y(\data_pdata[19]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3151));
 sg13g2_dfrbpq_1 \data_pdata[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3202),
    .D(net755),
    .Q(\data_pdata[19] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_mux2_1 \data_pdata[19]_sg13g2_mux2_1_A0  (.A0(\data_pdata[19] ),
    .A1(\data_pdata[27] ),
    .S(net3158),
    .X(\data_pdata[19]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_1 \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3149),
    .A2(\data_pdata[19]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\data_pdata[3]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_nand3b_1 \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C  (.B(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .C(\data_pdata[19]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ),
    .A_N(net3150));
 sg13g2_nand2_1 \data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B  (.Y(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .A(net2681),
    .B(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ));
 sg13g2_mux2_1 \data_pdata[19]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[19] ),
    .A1(net754),
    .S(net3049),
    .X(\data_pdata[19]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \data_pdata[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(net735),
    .Q(\data_pdata[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_mux2_1 \data_pdata[1]_sg13g2_mux2_1_A0  (.A0(\data_pdata[1] ),
    .A1(\data_pdata[9] ),
    .S(net3157),
    .X(\data_pdata[1]_sg13g2_mux2_1_A0_X ));
 sg13g2_nor2_1 \data_pdata[1]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B  (.A(net3149),
    .B(\data_pdata[1]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[1]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_mux2_1 \data_pdata[1]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[1] ),
    .A1(net734),
    .S(net3048),
    .X(\data_pdata[1]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \data_pdata[20]_sg13g2_a21oi_1_A2  (.A1(net3160),
    .A2(\data_pdata[20] ),
    .Y(\data_pdata[20]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3153));
 sg13g2_dfrbpq_1 \data_pdata[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(\data_pdata[20]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\data_pdata[20] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[20]_sg13g2_mux2_1_A0  (.A0(\data_pdata[20] ),
    .A1(\data_pdata[28] ),
    .S(net3160),
    .X(\data_pdata[20]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_2 \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2  (.B1(\data_pdata[4]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ),
    .Y(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[20]_sg13g2_mux2_1_A0_X ),
    .A1(net3153));
 sg13g2_nand3b_1 \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C  (.B(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .C(\data_pdata[20]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ),
    .A_N(net3152));
 sg13g2_nand2_2 \data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B  (.Y(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .A(net2683),
    .B(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y ));
 sg13g2_mux2_1 \data_pdata[20]_sg13g2_mux2_1_A1  (.A0(net907),
    .A1(net925),
    .S(net3050),
    .X(\data_pdata[20]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \data_pdata[21]_sg13g2_a21oi_1_A2  (.A1(net3155),
    .A2(\data_pdata[21] ),
    .Y(\data_pdata[21]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3150));
 sg13g2_dfrbpq_1 \data_pdata[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(net804),
    .Q(\data_pdata[21] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_mux2_1 \data_pdata[21]_sg13g2_mux2_1_A0  (.A0(\data_pdata[21] ),
    .A1(\data_pdata[29] ),
    .S(net3155),
    .X(\data_pdata[21]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_2 \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2  (.B1(\data_pdata[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ),
    .Y(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[21]_sg13g2_mux2_1_A0_X ),
    .A1(net3151));
 sg13g2_inv_1 \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A  (.Y(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y ),
    .A(\data_pdata[21]_sg13g2_mux2_1_A0_X ));
 sg13g2_o21ai_1 \data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2682),
    .Y(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y ),
    .A2(net3068));
 sg13g2_mux2_1 \data_pdata[21]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[21] ),
    .A1(net803),
    .S(net3049),
    .X(\data_pdata[21]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \data_pdata[22]_sg13g2_a21oi_1_A2  (.A1(net3162),
    .A2(\data_pdata[22] ),
    .Y(\data_pdata[22]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3154));
 sg13g2_dfrbpq_1 \data_pdata[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3204),
    .D(net799),
    .Q(\data_pdata[22] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[22]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[22] ),
    .A1(net798),
    .S(net3050),
    .X(\data_pdata[22]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2b_1 \data_pdata[22]_sg13g2_nor2b_1_B_N  (.A(net3162),
    .B_N(\data_pdata[22] ),
    .Y(\data_pdata[22]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_1 \data_pdata[23]_sg13g2_a21oi_1_A2  (.A1(net3160),
    .A2(\data_pdata[23] ),
    .Y(\data_pdata[23]_sg13g2_a21oi_1_A2_Y ),
    .B1(net3152));
 sg13g2_dfrbpq_1 \data_pdata[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net722),
    .Q(\data_pdata[23] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[23]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[23] ),
    .A1(net721),
    .S(net3050),
    .X(\data_pdata[23]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2b_1 \data_pdata[23]_sg13g2_nor2b_1_B_N  (.A(net3160),
    .B_N(\data_pdata[23] ),
    .Y(\data_pdata[23]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_2 \data_pdata[24]_sg13g2_a21oi_1_A2  (.B1(\data_pdata[16]_sg13g2_nor2b_1_B_N_Y ),
    .Y(\data_pdata[24]_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[24] ),
    .A1(net3159));
 sg13g2_a21oi_2 \data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2  (.B1(\data_pdata[0]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[24]_sg13g2_a21oi_1_A2_Y ),
    .A1(net3152));
 sg13g2_o21ai_1 \data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[24]_sg13g2_a21oi_1_A2_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_2 \data_pdata[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net928),
    .Q(\data_pdata[24] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[24]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[24] ),
    .A1(net927),
    .S(net3051),
    .X(\data_pdata[24]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[24]_sg13g2_nand2b_1_B  (.Y(\data_pdata[24]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[24] ),
    .A_N(net3159));
 sg13g2_o21ai_1 \data_pdata[24]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2683),
    .Y(\data_pdata[24]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[24]_sg13g2_nand2b_1_B_Y ),
    .A2(net3069));
 sg13g2_a21oi_1 \data_pdata[25]_sg13g2_a21oi_1_A2  (.A1(net3155),
    .A2(\data_pdata[25] ),
    .Y(\data_pdata[25]_sg13g2_a21oi_1_A2_Y ),
    .B1(\data_pdata[17]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_2 \data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2  (.B1(\data_pdata[1]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[25]_sg13g2_a21oi_1_A2_Y ),
    .A1(net3149));
 sg13g2_o21ai_1 \data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1  (.B1(net2682),
    .Y(\data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[25]_sg13g2_a21oi_1_A2_Y ),
    .A2(net3069));
 sg13g2_dfrbpq_2 \data_pdata[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net946),
    .Q(\data_pdata[25] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[25]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[25] ),
    .A1(net945),
    .S(net3048),
    .X(\data_pdata[25]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_2 \data_pdata[25]_sg13g2_nand2b_1_B  (.Y(\data_pdata[25]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[25] ),
    .A_N(net3155));
 sg13g2_o21ai_1 \data_pdata[25]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[25]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[25]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_1 \data_pdata[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net819),
    .Q(\data_pdata[26] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[26]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[26] ),
    .A1(net818),
    .S(net3048),
    .X(\data_pdata[26]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[26]_sg13g2_nand2b_1_B  (.Y(\data_pdata[26]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[26] ),
    .A_N(net3156));
 sg13g2_o21ai_1 \data_pdata[26]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[26]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[26]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_2 \data_pdata[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net942),
    .Q(\data_pdata[27] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_mux2_1 \data_pdata[27]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[27] ),
    .A1(net941),
    .S(net3049),
    .X(\data_pdata[27]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_2 \data_pdata[27]_sg13g2_nand2b_1_B  (.Y(\data_pdata[27]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[27] ),
    .A_N(net3158));
 sg13g2_o21ai_1 \data_pdata[27]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[27]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[27]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_2 \data_pdata[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3236),
    .D(\data_pdata[28]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\data_pdata[28] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[28]_sg13g2_mux2_1_A1  (.A0(net1051),
    .A1(net1083),
    .S(net3050),
    .X(\data_pdata[28]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_2 \data_pdata[28]_sg13g2_nand2b_1_B  (.Y(\data_pdata[28]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[28] ),
    .A_N(net3159));
 sg13g2_o21ai_1 \data_pdata[28]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[28]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[28]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_1 \data_pdata[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(net847),
    .Q(\data_pdata[29] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_mux2_1 \data_pdata[29]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[29] ),
    .A1(net846),
    .S(net3049),
    .X(\data_pdata[29]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[29]_sg13g2_nand2b_1_B  (.Y(\data_pdata[29]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[29] ),
    .A_N(net3155));
 sg13g2_o21ai_1 \data_pdata[29]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2682),
    .Y(\data_pdata[29]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[29]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_dfrbpq_1 \data_pdata[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3202),
    .D(net687),
    .Q(\data_pdata[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[2]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[2] ),
    .A1(net686),
    .S(net3048),
    .X(\data_pdata[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \data_pdata[2]_sg13g2_nor2_1_B  (.A(net3157),
    .B(\data_pdata[2] ),
    .Y(\data_pdata[2]_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \data_pdata[2]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C  (.A(net3149),
    .B(\data_pdata[10]_sg13g2_nor2b_1_A_Y ),
    .C(\data_pdata[2]_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[2]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_1 \data_pdata[30]_sg13g2_a21oi_1_A2  (.A1(net3162),
    .A2(\data_pdata[30] ),
    .Y(\data_pdata[30]_sg13g2_a21oi_1_A2_Y ),
    .B1(\data_pdata[22]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_2 \data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2  (.B1(\data_pdata[6]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[30]_sg13g2_a21oi_1_A2_Y ),
    .A1(net3154));
 sg13g2_o21ai_1 \data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1  (.B1(net2683),
    .Y(\data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[30]_sg13g2_a21oi_1_A2_Y ),
    .A2(net3069));
 sg13g2_dfrbpq_1 \data_pdata[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3204),
    .D(net1055),
    .Q(\data_pdata[30] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[30]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[30] ),
    .A1(net1054),
    .S(net3050),
    .X(\data_pdata[30]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_2 \data_pdata[30]_sg13g2_nand2b_1_B  (.Y(\data_pdata[30]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[30] ),
    .A_N(net3162));
 sg13g2_o21ai_1 \data_pdata[30]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2681),
    .Y(\data_pdata[30]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[30]_sg13g2_nand2b_1_B_Y ),
    .A2(net3068));
 sg13g2_a21oi_1 \data_pdata[31]_sg13g2_a21oi_1_A2  (.A1(net3160),
    .A2(\data_pdata[31] ),
    .Y(\data_pdata[31]_sg13g2_a21oi_1_A2_Y ),
    .B1(\data_pdata[23]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_2 \data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2  (.B1(\data_pdata[7]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[31]_sg13g2_a21oi_1_A2_Y ),
    .A1(net3152));
 sg13g2_o21ai_1 \data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1  (.B1(net2683),
    .Y(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[31]_sg13g2_a21oi_1_A2_Y ),
    .A2(net3069));
 sg13g2_dfrbpq_1 \data_pdata[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3233),
    .D(net859),
    .Q(\data_pdata[31] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_mux2_1 \data_pdata[31]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[31] ),
    .A1(net858),
    .S(net3050),
    .X(\data_pdata[31]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[31]_sg13g2_nand2b_1_B  (.Y(\data_pdata[31]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[31] ),
    .A_N(net3159));
 sg13g2_o21ai_1 \data_pdata[31]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1  (.B1(net2683),
    .Y(\data_pdata[31]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\data_pdata[31]_sg13g2_nand2b_1_B_Y ),
    .A2(net3069));
 sg13g2_dfrbpq_1 \data_pdata[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3202),
    .D(net689),
    .Q(\data_pdata[3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[3]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[3] ),
    .A1(net688),
    .S(net3048),
    .X(\data_pdata[3]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \data_pdata[3]_sg13g2_nor2_1_B  (.A(net3157),
    .B(\data_pdata[3] ),
    .Y(\data_pdata[3]_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \data_pdata[3]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C  (.A(net3149),
    .B(\data_pdata[11]_sg13g2_nor2b_1_A_Y ),
    .C(\data_pdata[3]_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[3]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_dfrbpq_1 \data_pdata[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(net699),
    .Q(\data_pdata[4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[4]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[4] ),
    .A1(net698),
    .S(net3051),
    .X(\data_pdata[4]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \data_pdata[4]_sg13g2_nor2_1_B  (.A(net3161),
    .B(\data_pdata[4] ),
    .Y(\data_pdata[4]_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \data_pdata[4]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C  (.A(net3153),
    .B(\data_pdata[12]_sg13g2_nor2b_1_A_Y ),
    .C(\data_pdata[4]_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[4]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_dfrbpq_1 \data_pdata[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net677),
    .Q(\data_pdata[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_mux2_1 \data_pdata[5]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[5] ),
    .A1(net676),
    .S(net3048),
    .X(\data_pdata[5]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \data_pdata[5]_sg13g2_nor2_1_B  (.A(net3157),
    .B(\data_pdata[5] ),
    .Y(\data_pdata[5]_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \data_pdata[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C  (.A(net3149),
    .B(\data_pdata[13]_sg13g2_nor2b_1_A_Y ),
    .C(\data_pdata[5]_sg13g2_nor2_1_B_Y ),
    .Y(\data_pdata[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_dfrbpq_1 \data_pdata[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(net720),
    .Q(\data_pdata[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_mux2_1 \data_pdata[6]_sg13g2_mux2_1_A0  (.A0(\data_pdata[6] ),
    .A1(\data_pdata[14] ),
    .S(net3162),
    .X(\data_pdata[6]_sg13g2_mux2_1_A0_X ));
 sg13g2_nor2_1 \data_pdata[6]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B  (.A(net3154),
    .B(\data_pdata[6]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[6]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_mux2_1 \data_pdata[6]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[6] ),
    .A1(net719),
    .S(net3051),
    .X(\data_pdata[6]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \data_pdata[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(net682),
    .Q(\data_pdata[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_mux2_1 \data_pdata[7]_sg13g2_mux2_1_A0  (.A0(\data_pdata[7] ),
    .A1(\data_pdata[15] ),
    .S(net3161),
    .X(\data_pdata[7]_sg13g2_mux2_1_A0_X ));
 sg13g2_nor2_1 \data_pdata[7]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B  (.A(net3153),
    .B(\data_pdata[7]_sg13g2_mux2_1_A0_X ),
    .Y(\data_pdata[7]_sg13g2_mux2_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_mux2_1 \data_pdata[7]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[7] ),
    .A1(net681),
    .S(net3051),
    .X(\data_pdata[7]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \data_pdata[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(net1148),
    .Q(\data_pdata[8] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_mux2_1 \data_pdata[8]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[8] ),
    .A1(net1147),
    .S(net3051),
    .X(\data_pdata[8]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[8]_sg13g2_nand2b_1_B  (.Y(\data_pdata[8]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[8] ),
    .A_N(net3159));
 sg13g2_a22oi_1 \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[24]_sg13g2_nand2b_1_B_Y ),
    .B2(net3152),
    .A2(\data_pdata[16]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[8]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21oi_2 \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.B1(net2714),
    .Y(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070));
 sg13g2_inv_2 \data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A  (.Y(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .A(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ));
 sg13g2_dfrbpq_1 \data_pdata[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3201),
    .D(net890),
    .Q(\data_pdata[9] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_mux2_1 \data_pdata[9]_sg13g2_mux2_1_A1  (.A0(\rsp_data_q[9] ),
    .A1(net889),
    .S(net3048),
    .X(\data_pdata[9]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \data_pdata[9]_sg13g2_nand2b_1_B  (.Y(\data_pdata[9]_sg13g2_nand2b_1_B_Y ),
    .B(\data_pdata[9] ),
    .A_N(net3157));
 sg13g2_a22oi_1 \data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\data_pdata[25]_sg13g2_nand2b_1_B_Y ),
    .B2(net3149),
    .A2(\data_pdata[17]_sg13g2_a21oi_1_A2_Y ),
    .A1(\data_pdata[9]_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21o_2 \data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2  (.A2(\data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y ),
    .A1(net3070),
    .B1(net2714),
    .X(\data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_dfrbpq_1 data_pvalid_sg13g2_dfrbpq_1_Q (.RESET_B(net3250),
    .D(data_pvalid_sg13g2_dfrbpq_1_Q_D),
    .Q(data_pvalid),
    .CLK(clknet_leaf_19_clk));
 sg13g2_inv_1 data_pvalid_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y (.Y(data_pvalid_sg13g2_dfrbpq_1_Q_D),
    .A(net3052));
 sg13g2_nand2b_2 data_pvalid_sg13g2_nand2b_1_B (.Y(data_pvalid_sg13g2_nand2b_1_B_Y),
    .B(net423),
    .A_N(\i_snitch.i_snitch_lsu.metadata_q[9] ));
 sg13g2_nor2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B (.A(\i_snitch.gpr_waddr[4] ),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y),
    .Y(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B (.A(net3163),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B (.A(\i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A_Y ),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X));
 sg13g2_nor3_2 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C (.A(net3163),
    .B(\i_snitch.gpr_waddr[4] ),
    .C(data_pvalid_sg13g2_nand2b_1_B_Y),
    .Y(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1_X));
 sg13g2_nor4_2 data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C (.A(net3163),
    .B(\i_snitch.gpr_waddr[4] ),
    .C(data_pvalid_sg13g2_nand2b_1_B_Y),
    .Y(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y),
    .D(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D));
 sg13g2_nor2_1 data_pvalid_sg13g2_nor2_1_A (.A(net423),
    .B(data_pvalid_sg13g2_nor2_1_A_B),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y));
 sg13g2_nor2_1 data_pvalid_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y (.A(net1408),
    .B(net2488),
    .Y(data_pvalid_sg13g2_nor2_1_A_B));
 sg13g2_dfrbpq_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D (.RESET_B(net3250),
    .D(data_pvalid_sg13g2_nor2_1_A_Y),
    .Q(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q),
    .CLK(clknet_leaf_20_clk));
 sg13g2_a21oi_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1 (.A1(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q),
    .A2(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_Y),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ));
 sg13g2_a221oi_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1 (.B2(net3141),
    .C1(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2),
    .B1(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_B1),
    .A1(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_and4_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .C(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .D(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D),
    .X(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1));
 sg13g2_nor2_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A_sg13g2_nor2_1_Y (.A(net3147),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A ),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A));
 sg13g2_nor3_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .C(net3007),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D));
 sg13g2_or2_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A_sg13g2_or2_1_X (.X(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A),
    .B(net3141),
    .A(net3144));
 sg13g2_nand2b_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B (.Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y),
    .B(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y),
    .A_N(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y ));
 sg13g2_or4_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B ),
    .B(net2719),
    .C(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_Y ),
    .D(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y),
    .X(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D_X));
 sg13g2_nand3_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1_Y ),
    .A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A_Y));
 sg13g2_nor2_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y (.A(net2848),
    .B(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2));
 sg13g2_nand3_1 data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y (.B(net2925),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ),
    .A(net2923),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B));
 sg13g2_nor2b_2 data_pvalid_sg13g2_nor2b_1_B_N (.A(\i_snitch.i_snitch_lsu.metadata_q[9] ),
    .B_N(data_pvalid),
    .Y(data_pvalid_sg13g2_nor2b_1_B_N_Y));
 sg13g2_and3_2 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C (.X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .A(net3163),
    .B(\i_snitch.gpr_waddr[4] ),
    .C(data_pvalid_sg13g2_nor2b_1_B_N_Y));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B (.A(\i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A_Y ),
    .B(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X));
 sg13g2_nand2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B (.Y(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y),
    .A(\i_snitch.gpr_waddr[4] ),
    .B(data_pvalid_sg13g2_nor2b_1_B_N_Y));
 sg13g2_nor2_2 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B (.A(net3163),
    .B(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y),
    .Y(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1_X));
 sg13g2_and2_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .B(\i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A_Y ),
    .X(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2_X));
 sg13g2_nor3_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B (.A(net3163),
    .B(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y),
    .C(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D),
    .Y(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B_Y));
 sg13g2_nand3_1 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C (.B(\i_snitch.gpr_waddr[4] ),
    .C(data_pvalid_sg13g2_nor2b_1_B_N_Y),
    .A(net3163),
    .Y(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y));
 sg13g2_nor2_2 data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D),
    .Y(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3245),
    .D(net748),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[0] ),
    .A1(net747),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(net1004),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[10] ),
    .A1(net1003),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(net874),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[11] ),
    .A1(net873),
    .S(net2914),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3245),
    .D(net1050),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[12] ),
    .A1(net1049),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(net1105),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[13] ),
    .A1(net1104),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3245),
    .D(net1090),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[14] ),
    .A1(net1089),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(net707),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[15] ),
    .A1(net706),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_nor2_1_B  (.A(net3177),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net950),
    .A1(net1069),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_nor2_1_B  (.A(net3174),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(net1043),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[17] ),
    .A1(net1042),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_nor2_1_B  (.A(net3175),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(net855),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[18] ),
    .A1(net854),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_nor2_1_B  (.A(net3175),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(net746),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[19] ),
    .A1(net745),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(net955),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[1] ),
    .A1(net954),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand3b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B_Y ),
    .A_N(net3178));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3248),
    .D(net1086),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net907),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3248),
    .D(net834),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[21] ),
    .A1(net833),
    .S(net2914),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(net1127),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[22] ),
    .A1(net1126),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(net837),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[23] ),
    .A1(net836),
    .S(net2914),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(net713),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[24] ),
    .A1(net712),
    .S(net2913),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(net1062),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[25] ),
    .A1(net1061),
    .S(net2916),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(net759),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[26] ),
    .A1(net758),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(net1066),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[27] ),
    .A1(net1065),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(net807),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[28] ),
    .A1(net806),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(net778),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[29] ),
    .A1(net777),
    .S(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(net961),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[2] ),
    .A1(net960),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(net776),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[30] ),
    .A1(net775),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(net832),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[31] ),
    .A1(net831),
    .S(net2917),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(net1140),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[3] ),
    .A1(net1139),
    .S(net2916),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(net1019),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[4] ),
    .A1(net1018),
    .S(net2916),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(net999),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[5] ),
    .A1(net998),
    .S(net2916),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3245),
    .D(net1134),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[6] ),
    .A1(net1133),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(net773),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[7] ),
    .A1(net772),
    .S(net2914),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(net771),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[8] ),
    .A1(net770),
    .S(net2915),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(net992),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\rsp_data_q[9] ),
    .A1(net991),
    .S(net2914),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_nor2_1_B  (.A(net3175),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_dfrbpq_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(net916),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ),
    .A(net915),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .A(net3177),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q ));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N  (.A(net3175),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_mux2_1_A1  (.A0(net747),
    .A1(net643),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A  (.B(net3178),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2 ),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_nand2_1_B_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B_Y ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2 ),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B_Y ));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1_sg13g2_or2_1_X  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B1 ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .A(net3179));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_B2 ),
    .B(net3179),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_B2 ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .A_N(net3178));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1_sg13g2_mux2_1_X  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ),
    .S(net3182),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_C1 ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B  (.A(net120),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B_X ));
 sg13g2_and3_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X ),
    .B(net2752),
    .A(net2849));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D  (.B(net2923),
    .C(net2926),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C  (.A(net3034),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A ),
    .D(net2922),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_and2_1_X  (.A(net116),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D  (.B(net3037),
    .C(net3073),
    .A(net3147),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B ));
 sg13g2_nor2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_nor2b_1_Y  (.A(net3147),
    .B_N(net3073),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A ));
 sg13g2_nor2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N  (.A(net2751),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net2848),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2 ),
    .A(net3073),
    .B(net2926));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B  (.A(net2848),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1 ),
    .B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_nand3b_1_B_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B1 ),
    .A(net3179),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_B2 ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .A_N(net3179));
 sg13g2_nand2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y ),
    .A(net114),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A ),
    .B(net3145),
    .A_N(net3142));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y ));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ),
    .B(net3141),
    .A_N(net3144));
 sg13g2_a22oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ),
    .B2(net2924),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_or2_1_X  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A ),
    .B(net3087),
    .A(net3085));
 sg13g2_or4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C_sg13g2_or4_1_X  (.A(net3083),
    .B(net3076),
    .C(net3079),
    .D(net3081),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ));
 sg13g2_a21o_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2  (.A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y ),
    .A1(net2815),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_or4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1 ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X ));
 sg13g2_nor4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C  (.A(net2710),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C_Y ));
 sg13g2_nor4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_D  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .B(net2744),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_or4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C  (.A(net2710),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2  (.B2(net2924),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1  (.B2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ),
    .C1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1 ),
    .A1(net2815),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net3148),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ));
 sg13g2_nor4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_D  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .B(net2744),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1_sg13g2_and4_1_X  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(net3035),
    .C(net3073),
    .D(net2926),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_B1 ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1_sg13g2_and4_1_X  (.A(net3035),
    .B(net2925),
    .C(net2922),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1 ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C  (.B(net2747),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_C ),
    .B(net3147),
    .A_N(net3142));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2 ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_A2 ),
    .A(net3034),
    .B(net2927));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1  (.A0(net1003),
    .A1(net576),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .S(net3177),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1  (.A0(net873),
    .A1(net655),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .S(net3177),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1049),
    .A1(net708),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .S(net118),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y ),
    .B(net118),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net3180),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ));
 sg13g2_and4_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and4_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(net3036),
    .C(net2927),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand4_1_A  (.B(net2927),
    .C(net3036),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_A ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1104),
    .A1(net822),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .S(net3180),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y ),
    .A(net3180),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1  (.B2(net3142),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ));
 sg13g2_nor4_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2 ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A ),
    .B(net3081),
    .A_N(net3075));
 sg13g2_or3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C  (.A(net3077),
    .B(net3079),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_Y ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C_sg13g2_nand3_1_Y  (.B(net3077),
    .C(net2927),
    .A(net3083),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_C ));
 sg13g2_or4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_or4_1_X  (.A(net3104),
    .B(net3125),
    .C(net3089),
    .D(net3093),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C_sg13g2_nand4_1_Y  (.B(net3083),
    .C(net3077),
    .A(net3085),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_C ),
    .D(net3079));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D_sg13g2_or2_1_X  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_D ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .A(net3087));
 sg13g2_or3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2 ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A_sg13g2_nand3_1_Y  (.B(net3073),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B ),
    .A(net3034),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A ));
 sg13g2_nand2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B ),
    .A(net3144),
    .B(net3141));
 sg13g2_nor3_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(net2750),
    .A_N(net86));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A  (.A(net86),
    .B_N(net2750),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .A_N(net3180));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1 ),
    .A1(net2923),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2 ));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2 ),
    .A2(net2924),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_A ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1 ),
    .A1(net96),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand4_1_Y  (.B(net2925),
    .C(net2922),
    .A(net3035),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_a21oi_1_A1_B1_sg13g2_o21ai_1_Y_B1 ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2 ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B ),
    .A(net3035),
    .B(net108));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B  (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_D_sg13g2_nor3_1_Y_A),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B_Y ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X  (.A(net3035),
    .B(net3141),
    .C(net108),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1 ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D_sg13g2_and2_1_X  (.A(net3147),
    .B(net3073),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_and4_1_X_D ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y ),
    .A(net3146),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1 ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_B ),
    .C(net98),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y  (.A(net96),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1 ));
 sg13g2_or4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B_sg13g2_or4_1_X  (.A(net3146),
    .B(net109),
    .C(net3085),
    .D(net3087),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B_sg13g2_nor2_1_Y  (.A(net2695),
    .B(net2748),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_B ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_and4_1_D  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1 ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C ));
 sg13g2_and3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A_sg13g2_and3_1_X  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A ),
    .A(net2924),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X ),
    .C(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_and2_1_X_A ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand3b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C  (.B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1 ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_B ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .A(net3034),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y  (.B(net2923),
    .C(net2926),
    .A(net3033),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A ),
    .D(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ));
 sg13g2_inv_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_inv_1_A  (.Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_B1),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2  (.B1(net2695),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1 ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_B_sg13g2_nor3_1_B_Y ),
    .A(net3141),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1 ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y  (.A(net3087),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y  (.B(net3079),
    .C(net3081),
    .A(net3085),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_A1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1  (.A0(net1089),
    .A1(net667),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .S(net3180),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1  (.A0(net706),
    .A1(net559),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3177),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1  (.A0(net1069),
    .A1(net552),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3174),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B  (.A(net3016),
    .B(net2997),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1  (.A0(net1042),
    .A1(net568),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3175),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_nor2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1  (.A0(net854),
    .A1(net561),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3175),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_nand2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A ),
    .A(net2963),
    .B(net2958));
 sg13g2_nand2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nand2_1_B_1  (.Y(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_B1 ),
    .A(net2972),
    .B(net2958));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_nor2_1_B  (.A(net2961),
    .B(net2954),
    .Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_B1 ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1  (.A0(net745),
    .A1(net564),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .S(net3177),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A_Y ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ),
    .B(net2720));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B  (.A(net2834),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ),
    .C(net2981),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B_sg13g2_nor2_1_Y  (.A(net3085),
    .B(net3087),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A  (.B(net2933),
    .C(net2919),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nand3_1_A_Y_sg13g2_o21ai_1_A2_B1 ),
    .A(net3083),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C_sg13g2_nor2_1_Y  (.A(net3083),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_C ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B_sg13g2_nand3_1_Y  (.B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ),
    .C(net2933),
    .A(net2941),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_A_B ));
 sg13g2_nor4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ),
    .C(net2810),
    .D(net2818),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y ),
    .A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y ));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ),
    .B(net92),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_and4_1_D  (.A(net3),
    .B(net1122),
    .C(net645),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ),
    .X(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B_Y ),
    .A(net645),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3245),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_mux2_1_A1  (.A0(net954),
    .A1(net605),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1409),
    .A1(net797),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .S(net3174),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3174),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .A2(net3174));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor2_1_B  (.A(net3107),
    .B(net2953),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_A2 ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net833),
    .A1(net702),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .S(net3176),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3176),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net3183),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1126),
    .A1(net1063),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .S(net3174),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3174),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net3174),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net836),
    .A1(net715),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .S(net3176),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_X ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A  (.A(net3088),
    .B(net3094),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2 ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3176),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net3176),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_B1 ),
    .A(net2930),
    .B(net2938));
 sg13g2_nand2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y ),
    .A(net2932),
    .B(net3096));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1  (.A0(net712),
    .A1(net622),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .S(net3177),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1  (.A0(net1061),
    .A1(net565),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .S(net3178),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1  (.A0(net758),
    .A1(net581),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .S(net3178),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1065),
    .A1(net697),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .S(net121),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y ),
    .B(net121),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net121),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ));
 sg13g2_nor4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ),
    .C(net51),
    .D(net2848),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_Y ));
 sg13g2_nor4_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_1  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_nor4_1_Y_A_sg13g2_or3_1_C_X ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .D(net2848));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1  (.A0(net806),
    .A1(net629),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .S(net3178),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1  (.A0(net777),
    .A1(net618),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .S(net3178),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3247),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net960),
    .A1(net751),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ),
    .S(net3180),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A  (.A(net114),
    .B(net3075),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_nand2_1_B_Y ),
    .A(net3179),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1  (.A0(net775),
    .A1(net608),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .S(net3181),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net831),
    .A1(net714),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .S(net121),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A  (.A(net3074),
    .B(net2537),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y ),
    .B(net121),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net121),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1139),
    .A1(net1093),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1  (.A0(net1018),
    .A1(net642),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ),
    .S(net3179),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3246),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1  (.A0(net998),
    .A1(net665),
    .S(net68),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .S(net3179),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2_1_A  (.A(net117),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A  (.A(net116),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1133),
    .A1(net869),
    .S(net2239),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .S(net118),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X_sg13g2_nor2_1_B  (.A(net3147),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ),
    .Y(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y ),
    .A(net3180),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .A_N(net3179));
 sg13g2_and4_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D  (.A(net3035),
    .B(net3147),
    .C(net2927),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X ));
 sg13g2_nand4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_nand4_1_D  (.B(net3036),
    .C(net2927),
    .A(net3147),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3242),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1  (.A0(net772),
    .A1(net586),
    .S(net2238),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .S(net3177),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1  (.A0(net770),
    .A1(net569),
    .S(net2240),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .S(net3178),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_mux2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1  (.A0(net991),
    .A1(net563),
    .S(net2237),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3176),
    .A_N(net563));
 sg13g2_nand2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_and2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .X(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2b_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_A ),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_and2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_and2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .X(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y_sg13g2_nor2_1_A  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ));
 sg13g2_dfrbpq_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ),
    .B(net125),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor2_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y  (.A(net3175),
    .B(net1319),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ));
 sg13g2_or3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X ));
 sg13g2_nor3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y  (.A(net2642),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2 ),
    .C1(net2957),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2962),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_mux4_1_X  (.S0(net3007),
    .A0(\i_snitch.sb_q[12] ),
    .A1(\i_snitch.sb_q[13] ),
    .A2(\i_snitch.sb_q[14] ),
    .A3(\i_snitch.sb_q[15] ),
    .S1(net2980),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(net3008));
 sg13g2_inv_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_snitch.sb_q[8] ));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.sb_q[9] ),
    .A2(net3008),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2980));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2 ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.sb_q[11] ),
    .B(net2803),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_A ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(net2969),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_nor2_1_Y_B ),
    .A1(\i_snitch.sb_q[10] ),
    .A2(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C ),
    .A1(net2837),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2_sg13g2_mux4_1_X  (.S0(net3007),
    .A0(\i_snitch.sb_q[4] ),
    .A1(\i_snitch.sb_q[5] ),
    .A2(\i_snitch.sb_q[6] ),
    .A3(\i_snitch.sb_q[7] ),
    .S1(net2980),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2832),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.sb_q[3] ),
    .B(net2803),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_a22oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(net2980),
    .B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .A2(net3008),
    .A1(\i_snitch.sb_q[1] ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_A_sg13g2_nor3_1_Y_C_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .B(net3032),
    .A_N(\i_snitch.sb_q[2] ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y  (.B2(net3089),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2634),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B ),
    .A2(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2939),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_mux4_1_X  (.S0(net3123),
    .A0(\i_snitch.sb_q[8] ),
    .A1(\i_snitch.sb_q[9] ),
    .A2(\i_snitch.sb_q[10] ),
    .A3(\i_snitch.sb_q[11] ),
    .S1(net3103),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a221oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .C1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A2(net2919));
 sg13g2_inv_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A1 ),
    .A(\i_snitch.sb_q[12] ));
 sg13g2_nand2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A(\i_snitch.sb_q[14] ),
    .B(net2949));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.sb_q[15] ),
    .A2(net3122),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .B1(net2941));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y  (.B1(net3093),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .A1(\i_snitch.sb_q[13] ),
    .A2(net2811));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1 ),
    .A1(net2818),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_mux4_1_X  (.S0(net3122),
    .A0(\i_snitch.sb_q[4] ),
    .A1(\i_snitch.sb_q[5] ),
    .A2(\i_snitch.sb_q[6] ),
    .A3(\i_snitch.sb_q[7] ),
    .S1(net3104),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.sb_q[2] ),
    .B(net3122),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_o21ai_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net3104),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A1(\i_snitch.sb_q[3] ),
    .A2(net2949));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.sb_q[1] ),
    .A2(net2826),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2823));
 sg13g2_a21o_2 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1  (.A2(net44),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ));
 sg13g2_and4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2 ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A ),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X  (.S0(net3072),
    .A0(\i_snitch.sb_q[12] ),
    .A1(\i_snitch.sb_q[13] ),
    .A2(\i_snitch.sb_q[14] ),
    .A3(\i_snitch.sb_q[15] ),
    .S1(net3071),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_A_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X  (.S0(net3072),
    .A0(\i_snitch.sb_q[8] ),
    .A1(\i_snitch.sb_q[9] ),
    .A2(\i_snitch.sb_q[10] ),
    .A3(\i_snitch.sb_q[11] ),
    .S1(net3071),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_B_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_nand2b_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .A_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_mux4_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N_sg13g2_mux4_1_X  (.S0(net3072),
    .A0(\i_snitch.sb_q[4] ),
    .A1(\i_snitch.sb_q[5] ),
    .A2(\i_snitch.sb_q[6] ),
    .A3(\i_snitch.sb_q[7] ),
    .S1(net3071),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_C_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y  (.A1(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2 ),
    .B1(net3072),
    .B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .A2(net3071),
    .A1(\i_snitch.sb_q[2] ));
 sg13g2_or2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_or2_1_X  (.X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .B(net3071),
    .A(\i_snitch.sb_q[1] ));
 sg13g2_nor2_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.sb_q[3] ),
    .B(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_A2_sg13g2_and4_1_X_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_B1  (.A1(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A_Y ),
    .A2(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B),
    .Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q_D ),
    .B1(net125));
 sg13g2_nand3_1 \i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A ),
    .C(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X ),
    .A(net78),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[37]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_snitch.pc_d[2] ),
    .Q(\i_req_arb.data_i[37] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_inv_2 \i_req_arb.data_i[37]_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ),
    .A(\i_req_arb.data_i[37] ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[38]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3261),
    .D(\i_snitch.pc_d[3] ),
    .Q(\i_req_arb.data_i[38] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[39]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3261),
    .D(\i_snitch.pc_d[4] ),
    .Q(\i_req_arb.data_i[39] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[40]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.pc_d[5] ),
    .Q(\i_req_arb.data_i[40] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_inv_2 \i_req_arb.data_i[40]_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .A(net1235));
 sg13g2_a21oi_1 \i_req_arb.data_i[41]_sg13g2_a21oi_1_B1  (.A1(net3086),
    .A2(net2536),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ),
    .B1(\i_req_arb.data_i[41] ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[41]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3257),
    .D(\i_snitch.pc_d[6] ),
    .Q(\i_req_arb.data_i[41] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_inv_2 \i_req_arb.data_i[41]_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ),
    .A(net1361));
 sg13g2_a221oi_1 \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1  (.B2(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2 ),
    .C1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1 ),
    .B1(net2637),
    .A1(\i_req_arb.data_i[42] ),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2721));
 sg13g2_a221oi_1 \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_o21ai_1_A1_Y ),
    .A1(net3089),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2 ),
    .A2(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A  (.Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y ),
    .A(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2 ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X ));
 sg13g2_inv_1 \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A  (.Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y ),
    .A(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y ));
 sg13g2_a21oi_1 \i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y  (.A1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ),
    .A2(net70),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[42]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_snitch.pc_d[7] ),
    .Q(\i_req_arb.data_i[42] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_inv_4 \i_req_arb.data_i[42]_sg13g2_inv_1_A  (.A(net1196),
    .Y(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[43]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3305),
    .D(\i_snitch.pc_d[8] ),
    .Q(\i_req_arb.data_i[43] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_a21o_1 \i_req_arb.data_i[44]_sg13g2_a21o_1_B1  (.A2(net100),
    .A1(net3080),
    .B1(\i_req_arb.data_i[44] ),
    .X(\i_req_arb.data_i[44]_sg13g2_a21o_1_B1_X ));
 sg13g2_dfrbpq_2 \i_req_arb.data_i[44]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.pc_d[9] ),
    .Q(\i_req_arb.data_i[44] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_nand3_1 \i_req_arb.data_i[44]_sg13g2_nand3_1_A  (.B(net3080),
    .C(net2537),
    .A(\i_req_arb.data_i[44] ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_a21o_2 \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X  (.A2(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ),
    .A1(net1331),
    .B1(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1 ),
    .X(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ));
 sg13g2_nor3_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y  (.A(net441),
    .B(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ),
    .C(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1 ));
 sg13g2_dfrbpq_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_inv_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A  (.Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_A_Y ),
    .A(net441));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y  (.A(net1392),
    .B(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B ),
    .Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net1332),
    .B(\i_req_arb.gen_arbiter.req_d[1] ),
    .Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B ));
 sg13g2_dfrbpq_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d ),
    .Q(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(net1332),
    .Q(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[1]_sg13g2_and2_1_B  (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ),
    .B(net1397),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_A ));
 sg13g2_dfrbpq_1 \i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(net1399),
    .Q(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_o21ai_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_o21ai_1_A2  (.B1(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ),
    .A2(\i_req_arb.gen_arbiter.req_d[1] ));
 sg13g2_or2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X  (.X(\i_req_arb.gen_arbiter.req_d[1] ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B ),
    .A(net1398));
 sg13g2_nor4_2 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y  (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_q ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B ),
    .D(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y ));
 sg13g2_a21o_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X  (.A2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2 ),
    .A1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1 ),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ));
 sg13g2_nand2b_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2 ),
    .A_N(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N ));
 sg13g2_nor3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A ));
 sg13g2_and3_2 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A  (.X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X ),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y ));
 sg13g2_nor2_2 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_nor2_1_Y  (.A(net2922),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B ));
 sg13g2_nand3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y ),
    .A(net44),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_Y ));
 sg13g2_inv_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B_sg13g2_inv_1_Y  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_B ),
    .A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nor2b_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A ),
    .B_N(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2 ));
 sg13g2_nand2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A ),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_nand3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B ),
    .C(net87),
    .A(net2928),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A ));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X  (.A(net3076),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B ),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B ));
 sg13g2_nand3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C  (.B(net3076),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_Y  (.A(net3079),
    .B(net3081),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B ));
 sg13g2_nand4_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C  (.B(net2924),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B ),
    .A(net2927),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_nand4_1_C_Y ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ));
 sg13g2_nor3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_or2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_or2_1_X  (.X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_B ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ));
 sg13g2_and3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C_sg13g2_and3_1_X  (.X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .A(net3076),
    .B(net3079),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y  (.B2(net2924),
    .C1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2744),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N ),
    .A2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand3b_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B ),
    .C(net2744),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B ),
    .A_N(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B_sg13g2_nand2_1_Y  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nand3b_1_A_N_B ),
    .A(net3076),
    .B(net3075));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2_sg13g2_nor2_1_Y  (.A(net3076),
    .B(net3075),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_and3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1_sg13g2_and3_1_X  (.X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B1 ),
    .A(net3033),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ));
 sg13g2_nor2b_2 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2_sg13g2_nor2b_1_Y  (.A(net3144),
    .B_N(net3142),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2 ));
 sg13g2_a21oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1  (.A1(net2744),
    .A2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_nand4_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C ),
    .A(net99),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y ),
    .D(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N ));
 sg13g2_and4_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C ),
    .D(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D ),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C ));
 sg13g2_nor2b_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N  (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N ),
    .B_N(net98),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_or2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D_sg13g2_or2_1_X  (.X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_D ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ),
    .A(net3141));
 sg13g2_nor3_2 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_nand4_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_A ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_C ),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B ),
    .D(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D ));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y ),
    .B(net2747),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_B ));
 sg13g2_a221oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D_sg13g2_a221oi_1_Y  (.B2(net2925),
    .C1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_A2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_B_Y ),
    .A1(net2922),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_D ),
    .A2(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ));
 sg13g2_a21oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1 ),
    .B1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net43),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1  (.B2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1 ),
    .C1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ),
    .A1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1 ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y ),
    .A2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2 ));
 sg13g2_nor3_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1_sg13g2_nor3_1_Y  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ),
    .C(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_B_Y_sg13g2_or4_1_D_X),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A1 ));
 sg13g2_inv_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2_sg13g2_inv_1_Y  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_A2 ),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B ));
 sg13g2_nand2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1_sg13g2_nand2_1_Y  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_B1 ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A  (.A(net44),
    .B(net2718),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1  (.Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_Y ),
    .B2(\i_req_arb.gen_arbiter.req_d[1] ),
    .A2(\i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2 ),
    .A1(net763));
 sg13g2_nand2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2_sg13g2_nand2_1_Y  (.Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_A2 ),
    .A(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ),
    .B(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ));
 sg13g2_dfrbpq_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3235),
    .D(\i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_arb.gen_arbiter.rr_q ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_inv_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_dfrbpq_1_Q_D ),
    .A(net764));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A  (.A(net763),
    .B(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B ),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_Y ));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B_sg13g2_and2_1_X  (.A(net1391),
    .B(net3172),
    .X(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_A  (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B ),
    .B(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ));
 sg13g2_o21ai_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1  (.B1(\i_req_arb.gen_arbiter.rr_q ),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B ),
    .A2(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_A ));
 sg13g2_a221oi_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2  (.B2(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ),
    .C1(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y ),
    .B1(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net3172));
 sg13g2_o21ai_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2  (.B1(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_Y),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1 ));
 sg13g2_inv_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1_sg13g2_inv_1_Y  (.Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1 ),
    .A(net2515));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .B(net42),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_or2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B  (.X(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B_X ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_and2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B  (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ),
    .B(net91),
    .X(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_2 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nand2_1_B  (.Y(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B),
    .A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ),
    .B(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_nor2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A  (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ),
    .B(net2496),
    .Y(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y ));
 sg13g2_or2_1 \i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A  (.X(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A_X ),
    .B(net2496),
    .A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_mux2_1 \i_req_register.data_o[38]_sg13g2_mux2_1_X  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38] ),
    .S(net3164),
    .X(\i_req_register.data_o[38] ));
 sg13g2_o21ai_1 \i_req_register.data_o[39]_sg13g2_o21ai_1_Y  (.B1(\i_req_register.data_o[39]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.data_o[39] ),
    .A1(net3173),
    .A2(\i_req_register.data_o[39]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_req_register.data_o[40]_sg13g2_mux2_1_X  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40] ),
    .S(net3165),
    .X(\i_req_register.data_o[40] ));
 sg13g2_o21ai_1 \i_req_register.data_o[41]_sg13g2_o21ai_1_Y  (.B1(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.data_o[41] ),
    .A1(net3164),
    .A2(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_req_register.data_o[42]_sg13g2_mux2_1_X  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42] ),
    .S(net3166),
    .X(\i_req_register.data_o[42] ));
 sg13g2_o21ai_1 \i_req_register.data_o[43]_sg13g2_o21ai_1_Y  (.B1(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.data_o[43] ),
    .A1(net3166),
    .A2(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.data_o[44]_sg13g2_o21ai_1_Y  (.B1(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.data_o[44] ),
    .A1(net3169),
    .A2(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.data_o[45]_sg13g2_o21ai_1_Y  (.B1(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.data_o[45] ),
    .A1(net3169),
    .A2(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_2 \i_req_register.data_o[5]_sg13g2_inv_1_A  (.Y(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ),
    .A(\i_req_register.data_o[5] ));
 sg13g2_nor2_2 \i_req_register.data_o[5]_sg13g2_inv_1_A_Y_sg13g2_nor2_1_B  (.A(net3053),
    .B(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ),
    .Y(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ));
 sg13g2_nor3_2 \i_req_register.data_o[5]_sg13g2_inv_1_A_Y_sg13g2_nor3_1_B  (.A(state),
    .B(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ),
    .C(req_data_valid_sg13g2_o21ai_1_Y_B1),
    .Y(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ));
 sg13g2_mux2_1 \i_req_register.data_o[5]_sg13g2_mux2_1_X  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .S(net3164),
    .X(\i_req_register.data_o[5] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_a21o_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21o_1_X  (.A2(net2491),
    .A1(net666),
    .B1(net2429),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2419),
    .A2(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2420));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2500),
    .B(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2482),
    .A2(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2532));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1263),
    .A2(net2494),
    .A1(net1193));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_and3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X  (.X(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ),
    .A(net2489),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2530),
    .A2(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2479));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net2429),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2489),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1365),
    .A2(net2491),
    .A1(net1258));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2422),
    .A2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2422));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2532),
    .A2(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2483));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1322),
    .A2(net2495),
    .A1(net1177));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B1(net2296),
    .B2(net1299),
    .A2(net2494),
    .A1(net1310));
 sg13g2_nand3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y  (.B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C ),
    .A(net2429),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y  (.B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B ),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C ),
    .A(net2490),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_B ),
    .A(net2500),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_Y_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .A1(net2481));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_C ),
    .A(net2421),
    .B(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3229),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2490),
    .A2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2481),
    .B(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2533),
    .C1(net2419),
    .B1(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .A1(net2500),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1183),
    .A2(net2494),
    .A1(net1156));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3188),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2489),
    .A2(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2530),
    .B(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2479),
    .C1(net2416),
    .B1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2499),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1343),
    .A2(net2491),
    .A1(net1377));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2417),
    .A2(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2417));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ),
    .B2(net2480),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ),
    .A1(net2498));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1336),
    .A2(net2492),
    .A1(net1287));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2417),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2417));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2531),
    .B(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ),
    .B2(net2480),
    .A2(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ),
    .A1(net2498));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1223),
    .A2(net2492),
    .A1(net1200));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2419),
    .A2(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2420));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2482),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .A1(net2532));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1306),
    .A2(net2494),
    .A1(net1240));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2416),
    .A2(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2415));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2479),
    .A2(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2530));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1388),
    .A2(net2491),
    .A1(net1283));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(net2489));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .A(net471),
    .B(net2491));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_o21ai_1_A2  (.B1(net3054),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ),
    .A1(net3167),
    .A2(net471));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2422),
    .A2(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2422));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2483),
    .A2(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2532));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2501),
    .B(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1297),
    .A2(net2495),
    .A1(net1187));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2421),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2421));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ),
    .B(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2481),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ),
    .A1(net2532));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1153),
    .A2(net2495),
    .A1(net1291));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2420),
    .A2(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2419));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2481),
    .A2(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ),
    .A1(net2533));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2502),
    .B(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net950),
    .A2(net2494),
    .A1(net1303));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3192),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2415),
    .A2(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2415));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2479),
    .A2(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2530));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1349),
    .A2(net2491),
    .A1(net1383));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2490),
    .A2(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2531),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2480),
    .C1(net2417),
    .B1(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ),
    .A1(net2498),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1226),
    .A2(net2495),
    .A1(net1233));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2418),
    .A2(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2418));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2480),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2498));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .B(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1362),
    .A2(net2492),
    .A1(net1207));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2490),
    .A2(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2481),
    .B(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2501),
    .C1(net2420),
    .B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2532),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net907),
    .A2(net2494),
    .A1(net1228));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2416),
    .A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2415));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2530),
    .A2(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2479));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1384),
    .A2(net2492),
    .A1(net1342));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2490),
    .A2(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2483),
    .B(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2501),
    .C1(net2422),
    .B1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2532),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1169),
    .A2(net2495),
    .A1(net1274));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2490),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y ));
 sg13g2_nor2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y  (.A(net2533),
    .B(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .B2(net2500),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ),
    .A1(net2481));
 sg13g2_nor2b_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_Y  (.A(net2490),
    .B_N(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1271),
    .A2(net2495),
    .A1(net1230));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3190),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net2429),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2493),
    .A1(net820));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1 ),
    .A(net2501));
 sg13g2_nor2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_and2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ),
    .A(net2501),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ));
 sg13g2_nand2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .A(net49),
    .B(net2515));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_o21ai_1_A2  (.B1(net3054),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ),
    .A1(net3168),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2420),
    .A2(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2419));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2500),
    .B(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .B2(net2533),
    .A2(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ),
    .A1(net2482));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1167),
    .A2(net2497),
    .A1(net1374));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2415),
    .A2(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2415));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2530),
    .A2(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2479));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1347),
    .A2(net2491),
    .A1(net1212));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2417),
    .A2(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2417));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2531),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ),
    .A1(net2480));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2498),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2298),
    .B2(net1330),
    .A2(net2495),
    .A1(net1217));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2417),
    .A2(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2418));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2531),
    .A2(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ),
    .A1(net2480));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2502),
    .B(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2295),
    .B2(net1345),
    .A2(net2492),
    .A1(net1265));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3229),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2426),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2419),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2419));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2532),
    .A2(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2481));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2500),
    .B(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2298),
    .B2(net1051),
    .A2(net2494),
    .A1(net1252));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_and3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X  (.X(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1 ),
    .A(net2489),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_B ),
    .A(net2499),
    .B(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ),
    .B2(net2479),
    .A2(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2530));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net2429),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2489),
    .A2(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1293),
    .A2(net2492),
    .A1(net1335));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2422),
    .A2(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2422));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2501),
    .A2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .A1(net2483));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .B(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2297),
    .B2(net1157),
    .A2(net2495),
    .A1(net1181));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2490),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2481),
    .C1(net2421),
    .B1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_nand2_1_A_Y_sg13g2_inv_1_A_Y ),
    .A1(net2500),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1107),
    .A2(net2497),
    .A1(net1269));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .C(net2429),
    .A(net2516),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2496),
    .B2(net1387),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ),
    .A1(net1378));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.data_o[39]_sg13g2_o21ai_1_Y_A2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2496),
    .A1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_inv_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ),
    .A(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2516),
    .A2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2427));
 sg13g2_inv_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_inv_1_A  (.Y(\i_req_register.data_o[39]_sg13g2_o21ai_1_Y_A2 ),
    .A(net1149));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_mux2_1_A0  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39] ),
    .A1(net579),
    .S(net2624),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3192),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2428),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2b_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .B_N(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A_sg13g2_nor2_1_Y  (.A(net49),
    .B(net2500),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .A(net537),
    .B(net2493));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_o21ai_1_A2  (.B1(net3054),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ),
    .A1(net3168),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_nor3_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2516),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ),
    .B1(net2427));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y  (.A(net1393),
    .B(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y  (.A(net1253),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_A2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2496),
    .A1(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2516),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2427));
 sg13g2_inv_4 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41]_sg13g2_inv_1_A  (.A(net931),
    .Y(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2429),
    .A1(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2b_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2_sg13g2_nand2b_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_B2 ),
    .B(net2516),
    .A_N(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(net1236),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_A2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2496),
    .A1(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2515),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2427));
 sg13g2_inv_4 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43]_sg13g2_inv_1_A  (.A(net844),
    .Y(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_A2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2497),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2516),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2427));
 sg13g2_inv_4 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44]_sg13g2_inv_1_A  (.A(net860),
    .Y(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3253),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_A2 ),
    .C1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2496),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_A1 ),
    .A(net1074));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2515),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2427));
 sg13g2_inv_4 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45]_sg13g2_inv_1_A  (.A(net768),
    .Y(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3190),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net2429),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2493),
    .A1(net533));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2 ),
    .A1(net2498),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y ),
    .B2(net94),
    .A2(net2496),
    .A1(net1380));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2425),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2420),
    .A2(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2419));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2502),
    .B(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2533),
    .A2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ),
    .A1(net2482));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2296),
    .B2(net1354),
    .A2(net2494),
    .A1(net1376));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2423),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2415),
    .A2(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(net2415));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2530),
    .B(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .B2(net2499),
    .A2(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(net2479));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1382),
    .A2(net2491),
    .A1(net1210));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2489),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2480),
    .B(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2498),
    .C1(net2418),
    .B1(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1369),
    .A2(net2492),
    .A1(net1208));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2424),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2489),
    .A2(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2480),
    .B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2498),
    .C1(net2418),
    .B1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_nor2b_1_Y_A ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2294),
    .B2(net1381),
    .A2(net2493),
    .A1(net1213));
 sg13g2_dfrbpq_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ),
    .A(net1392),
    .B(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nand2_1_A  (.Y(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ),
    .A(net1391),
    .B(net3172));
 sg13g2_nor2_2 \i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2_1_A  (.A(net1391),
    .B(net3164),
    .Y(req_data_valid_sg13g2_o21ai_1_Y_B1));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2  (.A1(net3165),
    .A2(net606),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_nor2b_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_B1_sg13g2_nor2b_1_Y  (.A(net3165),
    .B_N(net666),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3185),
    .D(net607),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .A1(net606),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(net578),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .A1(net577),
    .S(net2623),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net572),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .A1(net571),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .S(net3164),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net617),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .A1(net616),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .S(net3169),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net631),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .A1(net630),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .S(net3166),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(net650),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .A1(net649),
    .S(net2623),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(net575),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .A1(net574),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ),
    .S(net3165),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net624),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .A1(net623),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ),
    .S(net3166),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(net648),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .A1(net647),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ),
    .S(net3166),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(net595),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .A1(net594),
    .S(net2623),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(net680),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .A1(net679),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .S(net3173),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3185),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3167),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y ),
    .Y(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B2 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_mux2_1_A1  (.A0(net471),
    .A1(net609),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net592),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .A1(net591),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .S(net3169),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net585),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .A1(net584),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .S(net3169),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(net636),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .A1(net635),
    .S(net2623),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3192),
    .D(net663),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .A1(net662),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .S(net3168),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net583),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .A1(net582),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .S(net3169),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3197),
    .D(net626),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .A1(net625),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .S(net3166),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(net654),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .A1(net653),
    .S(net2624),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(net588),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .A1(net587),
    .S(net2618),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .S(net3168),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net611),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .A1(net610),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .S(net3170),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net604),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .A1(net603),
    .S(net2621),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .S(net3170),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3190),
    .D(net621),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3168),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y ),
    .Y(\strb_reg_q[2]_sg13g2_a21oi_1_A1_B1 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .A1(net620),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(net640),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .A1(net639),
    .S(net2624),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .S(net3171),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(net638),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .A1(net637),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .S(net3165),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(net599),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32] ),
    .A1(net598),
    .S(net2622),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32] ),
    .S(net3173),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net659),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33] ),
    .A1(net658),
    .S(net2622),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33] ),
    .S(net3170),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(net435),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y ),
    .A2(net2623),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34] ),
    .B(net2623),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y ),
    .A(net434));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3172),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(state));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(net437),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y ),
    .A2(net2618),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35] ),
    .B(net2618),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y ),
    .A(net436));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3165),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(state));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(net433),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y ),
    .A2(net2622),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36] ),
    .B(net2622),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y ),
    .A(net432));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3172),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(state));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3228),
    .D(net440),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y ),
    .A2(net2622),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37] ),
    .B(net2622),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y ),
    .A(net439));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3170),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(state));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net567),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38] ),
    .A1(net566),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(net580),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39]_sg13g2_nand2_1_B  (.Y(\i_req_register.data_o[39]_sg13g2_o21ai_1_Y_B1 ),
    .A(net3173),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3190),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y ),
    .A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3168),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y ),
    .Y(\strb_reg_q[4]_sg13g2_a21oi_1_A1_B1 ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_mux2_1_A1  (.A0(net537),
    .A1(net619),
    .S(net2617),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net628),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40] ),
    .A1(net627),
    .S(net2618),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net429),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_nand2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_A2 ),
    .A2(net2616));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_nand2_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_nand2_1_A_Y ),
    .A(net428),
    .B(net2616));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_nand2_1_B  (.Y(\i_req_register.data_o[41]_sg13g2_o21ai_1_Y_B1 ),
    .A(net3164),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net661),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42] ),
    .A1(net660),
    .S(net2620),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net425),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_nand2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_A2 ),
    .A2(net2619));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_nand2_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_nand2_1_A_Y ),
    .A(net424),
    .B(net2620));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_nand2_1_B  (.Y(\i_req_register.data_o[43]_sg13g2_o21ai_1_Y_B1 ),
    .A(net3166),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3200),
    .D(net431),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_nand2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_A2 ),
    .A2(net2621));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_nand2_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_nand2_1_A_Y ),
    .A(net430),
    .B(net2621));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_nand2_1_B  (.Y(\i_req_register.data_o[44]_sg13g2_o21ai_1_Y_B1 ),
    .A(net3169),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(net427),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_nand2_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_dfrbpq_1_Q_D ),
    .A1(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_A2 ),
    .A2(net2623));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_nand2_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_nand2_1_A_Y ),
    .A(net426),
    .B(net2623));
 sg13g2_nand2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_nand2_1_B  (.Y(\i_req_register.data_o[45]_sg13g2_o21ai_1_Y_B1 ),
    .A(net3169),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45] ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net446),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y ),
    .A2(net2617),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .B(net2617),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A  (.Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y ),
    .A(net445));
 sg13g2_a21oi_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2  (.A1(net3168),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y ),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(state));
 sg13g2_o21ai_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_B1  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .A1(net3168),
    .A2(net533));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(net590),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .A1(net589),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net613),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .A1(net612),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .S(net3166),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3188),
    .D(net602),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .A1(net601),
    .S(net2616),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .S(net3164),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(net652),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .A1(net651),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .S(net3167),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3196),
    .D(net633),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .A1(net632),
    .S(net2619),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_mux2_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1_1  (.A0(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .A1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ),
    .S(net3167),
    .X(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_dfrbpq_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3185),
    .D(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_nor2b_1 \i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2b_1_Y  (.A(req_data_valid_sg13g2_o21ai_1_Y_B1),
    .B_N(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B),
    .Y(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a22oi_1 \i_snitch.consec_pc[0]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.consec_pc[0]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2628),
    .B2(net49),
    .A2(net2755),
    .A1(\i_snitch.consec_pc[0] ));
 sg13g2_dfrbpq_2 \i_snitch.consec_pc[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3260),
    .D(\i_snitch.pc_d[0] ),
    .Q(\i_snitch.consec_pc[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3251),
    .D(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.gpr_waddr[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_a21oi_1 \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2487),
    .Y(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_2 \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .A(net3072));
 sg13g2_nor2_2 \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B  (.A(net3071),
    .B(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_1 \i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net1245),
    .B(net2487),
    .Y(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_dfrbpq_1 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3251),
    .D(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.gpr_waddr[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_a21oi_1 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2487),
    .Y(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_2 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .A(net3071));
 sg13g2_nor2_2 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A  (.A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_2 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1  (.A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1 ),
    .B(net3072),
    .Y(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ));
 sg13g2_nand2_2 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net3163),
    .B(net2487),
    .Y(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_dfrbpq_2 \i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3251),
    .D(\i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.gpr_waddr[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_a21oi_1 \i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .A2(net2488),
    .Y(\i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net1367),
    .B(net2488),
    .Y(\i_snitch.gpr_waddr[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2b_2 \i_snitch.gpr_waddr[6]_sg13g2_nor2b_1_A  (.A(\i_snitch.gpr_waddr[6] ),
    .B_N(\i_snitch.gpr_waddr[7] ),
    .Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_dfrbpq_2 \i_snitch.gpr_waddr[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3251),
    .D(\i_snitch.gpr_waddr[7]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.gpr_waddr[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_mux2_1 \i_snitch.gpr_waddr[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(net1389),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .S(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y ),
    .X(\i_snitch.gpr_waddr[7]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nand2_2 \i_snitch.gpr_waddr[7]_sg13g2_nand2_1_A  (.Y(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D),
    .A(\i_snitch.gpr_waddr[7] ),
    .B(\i_snitch.gpr_waddr[6] ));
 sg13g2_nor2_2 \i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A  (.A(\i_snitch.gpr_waddr[7] ),
    .B(\i_snitch.gpr_waddr[6] ),
    .Y(\i_snitch.gpr_waddr[7]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2b_2 \i_snitch.gpr_waddr[7]_sg13g2_nor2b_1_A  (.A(\i_snitch.gpr_waddr[7] ),
    .B_N(\i_snitch.gpr_waddr[6] ),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.i_snitch_lsu.handshake_pending_d ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A_sg13g2_nand2b_1_Y  (.Y(\i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A ),
    .B(net2515),
    .A_N(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_nor2_1_A_B ),
    .B(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_B ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_dfrbpq_1_Q  (.RESET_B(net3252),
    .D(\i_snitch.i_snitch_lsu.handshake_pending_d ),
    .Q(\i_snitch.i_snitch_lsu.handshake_pending_q ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_nor2_2 \i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A  (.A(net1407),
    .B(\i_snitch.i_snitch_lsu.handshake_pending_d_sg13g2_nor2_1_Y_A ),
    .Y(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2b_1 \i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A  (.A(net1407),
    .B_N(net1410),
    .Y(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2b_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_a21oi_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_X ),
    .A2(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand4_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A  (.B(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_B ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4] ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[0] ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y ),
    .D(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y ));
 sg13g2_inv_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_B_sg13g2_inv_1_Y  (.Y(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_B ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[1] ));
 sg13g2_nor2b_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .B_N(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nor2_1_A  (.A(net554),
    .B(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_or2_1 \i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_or2_1_A  (.X(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_or2_1_A_X ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[0] ));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_a21oi_1 \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ),
    .A2(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net1256),
    .B(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_nand2b_1_B  (.Y(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .A_N(net3151));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3204),
    .D(\i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_a21oi_1 \i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2531),
    .A2(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net3162),
    .B(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3204),
    .D(\i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_a21oi_1 \i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2486),
    .A2(net2501),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net3154),
    .B(net2486),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_inv_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_nand2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4] ),
    .B(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_or2_1_A_X ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .A1(net1160),
    .A2(net2488));
 sg13g2_nand3_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1 ));
 sg13g2_nand2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_C1 ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A ));
 sg13g2_nand4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y  (.B(net2925),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ),
    .A(net3034),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D ));
 sg13g2_xor2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D_sg13g2_xor2_1_X  (.B(net3141),
    .A(net3144),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A_sg13g2_nand4_1_Y_D ));
 sg13g2_nand3_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B  (.B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_B_A ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y ));
 sg13g2_nor4_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y ));
 sg13g2_and4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X  (.A(net2928),
    .B(net2924),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B ));
 sg13g2_and4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X  (.A(net3033),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D_sg13g2_nor2_1_Y  (.A(net3085),
    .B(net3083),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D_sg13g2_and4_1_X_D ));
 sg13g2_inv_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_inv_1_A  (.Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_A ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B ));
 sg13g2_and3_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X  (.X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C ),
    .A(net2923),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ));
 sg13g2_nor4_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B_sg13g2_nor4_1_Y  (.A(net3076),
    .B(net3080),
    .C(net3081),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ),
    .D(net3075));
 sg13g2_or2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B  (.X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A ));
 sg13g2_a21o_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1  (.A2(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2 ),
    .A1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1  (.Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2 ),
    .B2(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_B_sg13g2_and4_1_X_D ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2815));
 sg13g2_and2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_and2_1_X  (.A(net2923),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_and3_1_X_B ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2 ));
 sg13g2_and2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .B(net2815),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A ));
 sg13g2_or4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D ));
 sg13g2_and3_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A_sg13g2_and3_1_X  (.X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ),
    .A(net3035),
    .B(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ));
 sg13g2_and4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B_sg13g2_and4_1_X  (.A(net3034),
    .B(net2924),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_B ));
 sg13g2_a21o_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1  (.A2(net2815),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y ),
    .A2(net2815),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ));
 sg13g2_and4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_and4_1_X  (.A(net3033),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ),
    .D(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C ));
 sg13g2_and4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D_sg13g2_and4_1_X  (.A(net3035),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ),
    .D(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_D ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y_sg13g2_a21oi_1_A2  (.B1(net2928),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ),
    .A2(net70),
    .A1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nand2_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ),
    .A(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ),
    .B(net70));
 sg13g2_nand4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X ),
    .C(net2923),
    .A(net3034),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C_sg13g2_nor2_1_Y  (.A(net3145),
    .B(net3142),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C ));
 sg13g2_and2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B  (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B ),
    .X(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_X ));
 sg13g2_and2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_and2_1_B  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_B_Y_sg13g2_and2_1_B_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A ),
    .X(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A ));
 sg13g2_nand4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y  (.B(net2925),
    .C(net2926),
    .A(net3033),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A ),
    .D(net2922));
 sg13g2_nor2b_2 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D_sg13g2_nor2b_1_Y  (.A(net3142),
    .B_N(net3145),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B ),
    .A2(net3073));
 sg13g2_inv_4 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y_sg13g2_inv_1_A  (.A(net94),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A ),
    .B(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A1(net3077),
    .A2(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A(net2927),
    .B(net2744));
 sg13g2_nand3_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C  (.B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_A ),
    .C(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ));
 sg13g2_nand4_1 \i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand4_1_Y  (.B(net2925),
    .C(net2922),
    .A(net3033),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .D(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_D ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3251),
    .D(\i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_lsu.metadata_q[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_a21oi_1 \i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2488),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_nor2_1_A  (.A(net692),
    .B(net2488),
    .Y(\i_snitch.i_snitch_lsu.metadata_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[100] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2476),
    .C1(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2448),
    .A1(net2867),
    .Y(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[100]_sg13g2_nor3_1_A  (.A(net1305),
    .B(net2867),
    .C(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[100]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[100] ),
    .A2(net2803));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[101] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2408),
    .C1(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2448),
    .A1(net2866),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2906));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[101] ),
    .B(net2947),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor3_1_A  (.A(net1353),
    .B(net2866),
    .C(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[101] ),
    .A2(net2800));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2411),
    .B2(net1072),
    .A2(net2900),
    .A1(net2870));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3280),
    .D(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[102] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2450));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[102] ),
    .B(net2997),
    .Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[102]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[102] ),
    .A2(net2950));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2448),
    .B2(net2285),
    .A2(net2409),
    .A1(net1295));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3215),
    .D(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[103] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2866),
    .B(net2898));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[103] ),
    .B(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[103]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[103] ),
    .A2(net2947));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2410),
    .B2(net849),
    .A2(net2643),
    .A1(net2869));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[104] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2413));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[104] ),
    .B(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[104]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[104] ),
    .A2(net2952));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[105]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2410),
    .B2(net736),
    .A2(net2685),
    .A1(net2869));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[105] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2413));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[105] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y ),
    .A2(net2982),
    .Y(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net3027));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y ),
    .B2(net2282),
    .A2(net2411),
    .A1(net1302));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[106] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2870),
    .B(net2693));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[106] ),
    .B(net2953),
    .Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[106] ),
    .A2(net2804));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2833),
    .C1(net2639),
    .B1(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2955),
    .Y(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[107]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net817),
    .A2(net2680),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[107] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2413));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[107] ),
    .B(net2997),
    .Y(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2410),
    .B2(net1015),
    .A2(net2692),
    .A1(net2869));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[108] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2413));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[108] ),
    .A2(net2808));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2832),
    .C1(net2642),
    .B1(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2955),
    .Y(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(net2723),
    .A1(net3148));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2411),
    .B2(net1007),
    .A2(net2690),
    .A1(net2870));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[109] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2450));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[109] ),
    .A2(net2804));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2833),
    .C1(net2639),
    .B1(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2954),
    .Y(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2411),
    .B2(net911),
    .A2(net2688),
    .A1(net2870));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[110] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2450));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[110] ),
    .B(net2997),
    .Y(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net843),
    .A2(net2678),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[111] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2413));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[111] ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[111]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[111] ),
    .A2(net2952));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3289),
    .D(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[112] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2450),
    .B2(net2262),
    .A2(net2667),
    .A1(net2870));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net478),
    .B(net2411));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[112] ),
    .B(net2997),
    .Y(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[113]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2411),
    .B2(net922),
    .A2(net2664),
    .A1(net2870));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[113] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2413));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[113] ),
    .B(net2997),
    .Y(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2450),
    .B2(net2273),
    .A2(net2411),
    .A1(net1273));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[114] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2870),
    .B(net2676));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[114] ),
    .A2(net2805));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2833),
    .C1(net2639),
    .B1(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2954),
    .Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(net2724),
    .A1(net2955));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2448),
    .B2(net2271),
    .A2(net2409),
    .A1(net1165));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[115] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2866),
    .B(net2674));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[115] ),
    .A2(net2802));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2831),
    .C1(net2638),
    .B1(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2954),
    .Y(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[116]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net1060),
    .A2(net2671),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[116] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2414));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[116] ),
    .B(net2806),
    .Y(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2833),
    .Y(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2449),
    .B2(net2269),
    .A2(net2409),
    .A1(net1204));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[117] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2868),
    .B(net2670));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[117] ),
    .B(net2948),
    .Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_1  (.A(\i_snitch.i_snitch_regfile.mem[117] ),
    .B(net2802),
    .Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[118]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net982),
    .A2(net2651),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3320),
    .D(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[118] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2414));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[118] ),
    .B(net2806),
    .Y(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2833),
    .Y(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[119]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net1059),
    .A2(net2648),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3323),
    .D(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[119] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2414));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[119] ),
    .B(net2806),
    .Y(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2833),
    .Y(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2412),
    .B2(net1088),
    .A2(net2665),
    .A1(net2871));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[120] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2414));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[120] ),
    .B(net2952),
    .Y(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_1  (.A(\i_snitch.i_snitch_regfile.mem[120] ),
    .B(net2807),
    .Y(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2448),
    .B2(net2267),
    .A2(net2409),
    .A1(net1172));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3215),
    .D(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[121] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2866),
    .B(net2662));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[121] ),
    .B(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2448),
    .B2(net2255),
    .A2(net2409),
    .A1(net1250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[122] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2866),
    .B(net2660));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[122] ),
    .B(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2448),
    .B2(net2253),
    .A2(net2409),
    .A1(net1234));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[123] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2867),
    .B(net2658));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[123] ),
    .B(net2800),
    .Y(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2449),
    .B2(net2247),
    .A2(net2409),
    .A1(net1201));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[124] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2868),
    .B(net2656));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[124] ),
    .B(net2950),
    .Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_1  (.A(\i_snitch.i_snitch_regfile.mem[124] ),
    .B(net2801),
    .Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2450),
    .B2(net2251),
    .A2(net2410),
    .A1(net1180));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[125] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2868),
    .B(net2654));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[125] ),
    .B(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2450),
    .B2(net2245),
    .A2(net2411),
    .A1(net1216));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[126] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2870),
    .B(net2650));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[126] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y ),
    .A2(net2985),
    .Y(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net3028));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[127]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2410),
    .B2(net728),
    .A2(net2646),
    .A1(net2869));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[127] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2413));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[127] ),
    .B(net2802),
    .Y(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2832),
    .Y(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2352),
    .B2(net741),
    .A2(net2903),
    .A1(net2887));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[128] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0  (.S0(net3122),
    .A0(\i_snitch.i_snitch_regfile.mem[128] ),
    .A1(\i_snitch.i_snitch_regfile.mem[160] ),
    .A2(\i_snitch.i_snitch_regfile.mem[192] ),
    .A3(\i_snitch.i_snitch_regfile.mem[224] ),
    .S1(net3104),
    .X(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1  (.S0(net3007),
    .A0(\i_snitch.i_snitch_regfile.mem[128] ),
    .A1(\i_snitch.i_snitch_regfile.mem[160] ),
    .A2(\i_snitch.i_snitch_regfile.mem[192] ),
    .A3(\i_snitch.i_snitch_regfile.mem[224] ),
    .S1(net2981),
    .X(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B  (.A(net2837),
    .B(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2818),
    .B(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[129] ),
    .A2(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y ),
    .B1(net3013));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y  (.A(net2971),
    .B(net2955),
    .Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_1_X ),
    .B2(net3107),
    .A2(net2920),
    .A1(\i_snitch.i_snitch_regfile.mem[129] ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_A2_sg13g2_nor2_1_Y  (.A(net3127),
    .B(net3106),
    .Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_A2 ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_nand2_1_A_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(net2817));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[129] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2446),
    .B2(net2513),
    .A2(net2901),
    .A1(net2888));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[129]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net463),
    .B(net2350));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[130] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2445),
    .A1(net2885),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0  (.S0(net3001),
    .A0(\i_snitch.i_snitch_regfile.mem[130] ),
    .A1(\i_snitch.i_snitch_regfile.mem[162] ),
    .A2(\i_snitch.i_snitch_regfile.mem[194] ),
    .A3(\i_snitch.i_snitch_regfile.mem[226] ),
    .S1(net2974),
    .X(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1  (.S0(net3117),
    .A0(\i_snitch.i_snitch_regfile.mem[130] ),
    .A1(\i_snitch.i_snitch_regfile.mem[162] ),
    .A2(\i_snitch.i_snitch_regfile.mem[194] ),
    .A3(\i_snitch.i_snitch_regfile.mem[226] ),
    .S1(net3099),
    .X(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net2962),
    .C1(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ),
    .A1(net3093),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2751));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[130]_sg13g2_nor3_1_A  (.A(net1286),
    .B(net2885),
    .C(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[131] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2447),
    .A1(net2886),
    .Y(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0  (.S0(net3006),
    .A0(\i_snitch.i_snitch_regfile.mem[131] ),
    .A1(\i_snitch.i_snitch_regfile.mem[163] ),
    .A2(\i_snitch.i_snitch_regfile.mem[195] ),
    .A3(\i_snitch.i_snitch_regfile.mem[227] ),
    .S1(net2979),
    .X(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1  (.S0(net3120),
    .A0(\i_snitch.i_snitch_regfile.mem[131] ),
    .A1(\i_snitch.i_snitch_regfile.mem[163] ),
    .A2(\i_snitch.i_snitch_regfile.mem[195] ),
    .A3(\i_snitch.i_snitch_regfile.mem[227] ),
    .S1(net3101),
    .X(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B  (.A(net2817),
    .B(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[131]_sg13g2_nor3_1_A  (.A(net1289),
    .B(net2886),
    .C(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[132] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2445),
    .A1(net2887),
    .Y(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0  (.S0(net3007),
    .A0(\i_snitch.i_snitch_regfile.mem[132] ),
    .A1(\i_snitch.i_snitch_regfile.mem[164] ),
    .A2(\i_snitch.i_snitch_regfile.mem[196] ),
    .A3(\i_snitch.i_snitch_regfile.mem[228] ),
    .S1(net2980),
    .X(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1  (.S0(net3122),
    .A0(\i_snitch.i_snitch_regfile.mem[132] ),
    .A1(\i_snitch.i_snitch_regfile.mem[164] ),
    .A2(\i_snitch.i_snitch_regfile.mem[196] ),
    .A3(\i_snitch.i_snitch_regfile.mem[228] ),
    .S1(net3104),
    .X(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2837),
    .A2(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[132]_sg13g2_nor3_1_A  (.A(net1247),
    .B(net2890),
    .C(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[133] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2445),
    .A1(net2885),
    .Y(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0  (.S0(net3117),
    .A0(\i_snitch.i_snitch_regfile.mem[133] ),
    .A1(\i_snitch.i_snitch_regfile.mem[165] ),
    .A2(\i_snitch.i_snitch_regfile.mem[197] ),
    .A3(\i_snitch.i_snitch_regfile.mem[229] ),
    .S1(net3099),
    .X(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1  (.S0(net3001),
    .A0(\i_snitch.i_snitch_regfile.mem[133] ),
    .A1(\i_snitch.i_snitch_regfile.mem[165] ),
    .A2(\i_snitch.i_snitch_regfile.mem[197] ),
    .A3(\i_snitch.i_snitch_regfile.mem[229] ),
    .S1(net2974),
    .X(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[101]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2816),
    .A2(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[133]_sg13g2_nor3_1_A  (.A(net1370),
    .B(net2885),
    .C(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2350),
    .B2(net965),
    .A2(net2900),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[134] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2446));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0  (.S0(net124),
    .A0(\i_snitch.i_snitch_regfile.mem[134] ),
    .A1(\i_snitch.i_snitch_regfile.mem[166] ),
    .A2(\i_snitch.i_snitch_regfile.mem[198] ),
    .A3(\i_snitch.i_snitch_regfile.mem[230] ),
    .S1(net3107),
    .X(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1  (.S0(net3013),
    .A0(\i_snitch.i_snitch_regfile.mem[134] ),
    .A1(\i_snitch.i_snitch_regfile.mem[166] ),
    .A2(\i_snitch.i_snitch_regfile.mem[198] ),
    .A3(\i_snitch.i_snitch_regfile.mem[230] ),
    .S1(net2986),
    .X(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net938),
    .A2(net2445),
    .A1(net2284));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3191),
    .D(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[135] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2886),
    .B(net2897));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[135] ),
    .A1(\i_snitch.i_snitch_regfile.mem[167] ),
    .A2(\i_snitch.i_snitch_regfile.mem[199] ),
    .A3(\i_snitch.i_snitch_regfile.mem[231] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1  (.S0(net2999),
    .A0(\i_snitch.i_snitch_regfile.mem[135] ),
    .A1(\i_snitch.i_snitch_regfile.mem[167] ),
    .A2(\i_snitch.i_snitch_regfile.mem[199] ),
    .A3(\i_snitch.i_snitch_regfile.mem[231] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[103]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_X ),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2352),
    .B2(net752),
    .A2(net2643),
    .A1(net2887));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[136] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0  (.S0(net3123),
    .A0(\i_snitch.i_snitch_regfile.mem[136] ),
    .A1(\i_snitch.i_snitch_regfile.mem[168] ),
    .A2(\i_snitch.i_snitch_regfile.mem[200] ),
    .A3(\i_snitch.i_snitch_regfile.mem[232] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1  (.S0(net3008),
    .A0(\i_snitch.i_snitch_regfile.mem[136] ),
    .A1(\i_snitch.i_snitch_regfile.mem[168] ),
    .A2(\i_snitch.i_snitch_regfile.mem[200] ),
    .A3(\i_snitch.i_snitch_regfile.mem[232] ),
    .S1(net2982),
    .X(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2837),
    .A2(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1  (.A2(net2753),
    .A1(net3081),
    .B1(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2818),
    .B(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2352),
    .B2(net738),
    .A2(net2686),
    .A1(net2887));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[137] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0  (.S0(net3124),
    .A0(\i_snitch.i_snitch_regfile.mem[137] ),
    .A1(\i_snitch.i_snitch_regfile.mem[169] ),
    .A2(\i_snitch.i_snitch_regfile.mem[201] ),
    .A3(\i_snitch.i_snitch_regfile.mem[233] ),
    .S1(net3103),
    .X(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1  (.S0(net3009),
    .A0(\i_snitch.i_snitch_regfile.mem[137] ),
    .A1(\i_snitch.i_snitch_regfile.mem[169] ),
    .A2(\i_snitch.i_snitch_regfile.mem[201] ),
    .A3(\i_snitch.i_snitch_regfile.mem[233] ),
    .S1(net2983),
    .X(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .A_N(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2818),
    .B(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net852),
    .A2(net2446),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3278),
    .D(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[138] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2889),
    .B(net2693));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0  (.S0(net3128),
    .A0(\i_snitch.i_snitch_regfile.mem[138] ),
    .A1(\i_snitch.i_snitch_regfile.mem[170] ),
    .A2(\i_snitch.i_snitch_regfile.mem[202] ),
    .A3(\i_snitch.i_snitch_regfile.mem[234] ),
    .S1(net3107),
    .X(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1  (.S0(net3014),
    .A0(\i_snitch.i_snitch_regfile.mem[138] ),
    .A1(\i_snitch.i_snitch_regfile.mem[170] ),
    .A2(\i_snitch.i_snitch_regfile.mem[202] ),
    .A3(\i_snitch.i_snitch_regfile.mem[234] ),
    .S1(net2986),
    .X(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ),
    .A(net3078),
    .B(net2753));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[106]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2819),
    .A2(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net1097),
    .A2(net2679),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[139] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0  (.S0(net3136),
    .A0(\i_snitch.i_snitch_regfile.mem[139] ),
    .A1(\i_snitch.i_snitch_regfile.mem[171] ),
    .A2(\i_snitch.i_snitch_regfile.mem[203] ),
    .A3(\i_snitch.i_snitch_regfile.mem[235] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1  (.S0(net3021),
    .A0(\i_snitch.i_snitch_regfile.mem[139] ),
    .A1(\i_snitch.i_snitch_regfile.mem[171] ),
    .A2(\i_snitch.i_snitch_regfile.mem[203] ),
    .A3(\i_snitch.i_snitch_regfile.mem[235] ),
    .S1(net2992),
    .X(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[107]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net740),
    .A2(net2692),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3310),
    .D(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[140] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0  (.S0(net3133),
    .A0(\i_snitch.i_snitch_regfile.mem[140] ),
    .A1(\i_snitch.i_snitch_regfile.mem[172] ),
    .A2(\i_snitch.i_snitch_regfile.mem[204] ),
    .A3(\i_snitch.i_snitch_regfile.mem[236] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1  (.S0(net3019),
    .A0(\i_snitch.i_snitch_regfile.mem[140] ),
    .A1(\i_snitch.i_snitch_regfile.mem[172] ),
    .A2(\i_snitch.i_snitch_regfile.mem[204] ),
    .A3(\i_snitch.i_snitch_regfile.mem[236] ),
    .S1(net2990),
    .X(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .A_N(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net959),
    .A2(net2689),
    .A1(net2889));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[141] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2446));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0  (.S0(net3130),
    .A0(\i_snitch.i_snitch_regfile.mem[141] ),
    .A1(\i_snitch.i_snitch_regfile.mem[173] ),
    .A2(\i_snitch.i_snitch_regfile.mem[205] ),
    .A3(\i_snitch.i_snitch_regfile.mem[237] ),
    .S1(net3108),
    .X(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1  (.S0(net3017),
    .A0(\i_snitch.i_snitch_regfile.mem[141] ),
    .A1(\i_snitch.i_snitch_regfile.mem[173] ),
    .A2(\i_snitch.i_snitch_regfile.mem[205] ),
    .A3(\i_snitch.i_snitch_regfile.mem[237] ),
    .S1(net2988),
    .X(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[109]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_A ),
    .A(net73),
    .B(net2724));
 sg13g2_inv_2 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net1116),
    .A2(net2688),
    .A1(net2889));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3289),
    .D(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[142] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2446));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0  (.S0(net3130),
    .A0(\i_snitch.i_snitch_regfile.mem[142] ),
    .A1(\i_snitch.i_snitch_regfile.mem[174] ),
    .A2(\i_snitch.i_snitch_regfile.mem[206] ),
    .A3(\i_snitch.i_snitch_regfile.mem[238] ),
    .S1(net3109),
    .X(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1  (.S0(net3018),
    .A0(\i_snitch.i_snitch_regfile.mem[142] ),
    .A1(\i_snitch.i_snitch_regfile.mem[174] ),
    .A2(\i_snitch.i_snitch_regfile.mem[206] ),
    .A3(\i_snitch.i_snitch_regfile.mem[238] ),
    .S1(net2989),
    .X(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[110]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2639),
    .B(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2725),
    .A1(net74));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2352),
    .B2(net1142),
    .A2(net2678),
    .A1(net2890));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3299),
    .D(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[143] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0  (.S0(net3136),
    .A0(\i_snitch.i_snitch_regfile.mem[143] ),
    .A1(\i_snitch.i_snitch_regfile.mem[175] ),
    .A2(\i_snitch.i_snitch_regfile.mem[207] ),
    .A3(\i_snitch.i_snitch_regfile.mem[239] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1  (.S0(net3021),
    .A0(\i_snitch.i_snitch_regfile.mem[143] ),
    .A1(\i_snitch.i_snitch_regfile.mem[175] ),
    .A2(\i_snitch.i_snitch_regfile.mem[207] ),
    .A3(\i_snitch.i_snitch_regfile.mem[239] ),
    .S1(net2992),
    .X(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1  (.A2(net2724),
    .A1(net3022),
    .B1(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net1047),
    .A2(net2446),
    .A1(net2262));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[144] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2889),
    .B(net2667));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0  (.S0(net3129),
    .A0(\i_snitch.i_snitch_regfile.mem[144] ),
    .A1(\i_snitch.i_snitch_regfile.mem[176] ),
    .A2(\i_snitch.i_snitch_regfile.mem[208] ),
    .A3(\i_snitch.i_snitch_regfile.mem[240] ),
    .S1(net3108),
    .X(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1  (.S0(net3016),
    .A0(\i_snitch.i_snitch_regfile.mem[144] ),
    .A1(\i_snitch.i_snitch_regfile.mem[176] ),
    .A2(\i_snitch.i_snitch_regfile.mem[208] ),
    .A3(\i_snitch.i_snitch_regfile.mem[240] ),
    .S1(net2987),
    .X(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[112]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2352),
    .B2(net767),
    .A2(net2663),
    .A1(net2890));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[145] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0  (.S0(net3136),
    .A0(\i_snitch.i_snitch_regfile.mem[145] ),
    .A1(\i_snitch.i_snitch_regfile.mem[177] ),
    .A2(\i_snitch.i_snitch_regfile.mem[209] ),
    .A3(\i_snitch.i_snitch_regfile.mem[241] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1  (.S0(net3021),
    .A0(\i_snitch.i_snitch_regfile.mem[145] ),
    .A1(\i_snitch.i_snitch_regfile.mem[177] ),
    .A2(\i_snitch.i_snitch_regfile.mem[209] ),
    .A3(\i_snitch.i_snitch_regfile.mem[241] ),
    .S1(net2994),
    .X(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[113]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2639),
    .B(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1  (.A2(net2724),
    .A1(net2965),
    .B1(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net828),
    .A2(net2447),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[146] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2889),
    .B(net2675));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0  (.S0(net3129),
    .A0(\i_snitch.i_snitch_regfile.mem[146] ),
    .A1(\i_snitch.i_snitch_regfile.mem[178] ),
    .A2(\i_snitch.i_snitch_regfile.mem[210] ),
    .A3(\i_snitch.i_snitch_regfile.mem[242] ),
    .S1(net3108),
    .X(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1  (.S0(net3016),
    .A0(\i_snitch.i_snitch_regfile.mem[146] ),
    .A1(\i_snitch.i_snitch_regfile.mem[178] ),
    .A2(\i_snitch.i_snitch_regfile.mem[210] ),
    .A3(\i_snitch.i_snitch_regfile.mem[242] ),
    .S1(net2987),
    .X(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .A_N(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[146]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net1033),
    .A2(net2445),
    .A1(net2270));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3190),
    .D(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[147] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2885),
    .B(net2673));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[147] ),
    .A1(\i_snitch.i_snitch_regfile.mem[179] ),
    .A2(\i_snitch.i_snitch_regfile.mem[211] ),
    .A3(\i_snitch.i_snitch_regfile.mem[243] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1  (.S0(net2999),
    .A0(\i_snitch.i_snitch_regfile.mem[147] ),
    .A1(\i_snitch.i_snitch_regfile.mem[179] ),
    .A2(\i_snitch.i_snitch_regfile.mem[211] ),
    .A3(\i_snitch.i_snitch_regfile.mem[243] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[115]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nand2_1_A_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net871),
    .A2(net2671),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[148] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2348));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0  (.S0(net3138),
    .A0(\i_snitch.i_snitch_regfile.mem[148] ),
    .A1(\i_snitch.i_snitch_regfile.mem[180] ),
    .A2(\i_snitch.i_snitch_regfile.mem[212] ),
    .A3(\i_snitch.i_snitch_regfile.mem[244] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1  (.S0(net3022),
    .A0(\i_snitch.i_snitch_regfile.mem[148] ),
    .A1(\i_snitch.i_snitch_regfile.mem[180] ),
    .A2(\i_snitch.i_snitch_regfile.mem[212] ),
    .A3(\i_snitch.i_snitch_regfile.mem[244] ),
    .S1(net2993),
    .X(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[116]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1  (.A1(net3134),
    .A2(net2849),
    .Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net1087),
    .A2(net2447),
    .A1(net2268));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[149] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2886),
    .B(net2669));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0  (.S0(net3119),
    .A0(\i_snitch.i_snitch_regfile.mem[149] ),
    .A1(\i_snitch.i_snitch_regfile.mem[181] ),
    .A2(\i_snitch.i_snitch_regfile.mem[213] ),
    .A3(\i_snitch.i_snitch_regfile.mem[245] ),
    .S1(net3101),
    .X(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1  (.S0(net3005),
    .A0(\i_snitch.i_snitch_regfile.mem[149] ),
    .A1(\i_snitch.i_snitch_regfile.mem[181] ),
    .A2(\i_snitch.i_snitch_regfile.mem[213] ),
    .A3(\i_snitch.i_snitch_regfile.mem[245] ),
    .S1(net2978),
    .X(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2837),
    .A2(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net3105),
    .C1(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2850),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2754));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2817),
    .A2(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net853),
    .A2(net2651),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[150] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2348));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0  (.S0(net3138),
    .A0(\i_snitch.i_snitch_regfile.mem[150] ),
    .A1(\i_snitch.i_snitch_regfile.mem[182] ),
    .A2(\i_snitch.i_snitch_regfile.mem[214] ),
    .A3(\i_snitch.i_snitch_regfile.mem[246] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1  (.S0(net3023),
    .A0(\i_snitch.i_snitch_regfile.mem[150] ),
    .A1(\i_snitch.i_snitch_regfile.mem[182] ),
    .A2(\i_snitch.i_snitch_regfile.mem[214] ),
    .A3(\i_snitch.i_snitch_regfile.mem[246] ),
    .S1(net2994),
    .X(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[118]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2849),
    .A1(net3096));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1 ),
    .B2(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2 ),
    .A2(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .C(net2548),
    .A(net2569),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a22oi_1_A2_B2 ),
    .A1(net2565),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net851),
    .A2(net2648),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[151] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2348));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0  (.S0(net3137),
    .A0(\i_snitch.i_snitch_regfile.mem[151] ),
    .A1(\i_snitch.i_snitch_regfile.mem[183] ),
    .A2(\i_snitch.i_snitch_regfile.mem[215] ),
    .A3(\i_snitch.i_snitch_regfile.mem[247] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1  (.S0(net3022),
    .A0(\i_snitch.i_snitch_regfile.mem[151] ),
    .A1(\i_snitch.i_snitch_regfile.mem[183] ),
    .A2(\i_snitch.i_snitch_regfile.mem[215] ),
    .A3(\i_snitch.i_snitch_regfile.mem[247] ),
    .S1(net2993),
    .X(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[119]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2820),
    .B(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2350),
    .B2(net732),
    .A2(net2665),
    .A1(net2888));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[152] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2348));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0  (.S0(net3137),
    .A0(\i_snitch.i_snitch_regfile.mem[152] ),
    .A1(\i_snitch.i_snitch_regfile.mem[184] ),
    .A2(\i_snitch.i_snitch_regfile.mem[216] ),
    .A3(\i_snitch.i_snitch_regfile.mem[248] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1  (.S0(net3022),
    .A0(\i_snitch.i_snitch_regfile.mem[152] ),
    .A1(\i_snitch.i_snitch_regfile.mem[184] ),
    .A2(\i_snitch.i_snitch_regfile.mem[216] ),
    .A3(\i_snitch.i_snitch_regfile.mem[248] ),
    .S1(net2993),
    .X(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2839),
    .A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .C1(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2849),
    .A1(net3074),
    .Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2753));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net1151),
    .A2(net2445),
    .A1(net2266));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[153] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2885),
    .B(net2661));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0  (.S0(net3116),
    .A0(\i_snitch.i_snitch_regfile.mem[153] ),
    .A1(\i_snitch.i_snitch_regfile.mem[185] ),
    .A2(\i_snitch.i_snitch_regfile.mem[217] ),
    .A3(\i_snitch.i_snitch_regfile.mem[249] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1  (.S0(net3000),
    .A0(\i_snitch.i_snitch_regfile.mem[153] ),
    .A1(\i_snitch.i_snitch_regfile.mem[185] ),
    .A2(\i_snitch.i_snitch_regfile.mem[217] ),
    .A3(\i_snitch.i_snitch_regfile.mem[249] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[121]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ),
    .C1(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2849),
    .A1(net3074),
    .Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2752));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net1009),
    .A2(net2445),
    .A1(net2254));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[154] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2885),
    .B(net2659));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[154] ),
    .A1(\i_snitch.i_snitch_regfile.mem[186] ),
    .A2(\i_snitch.i_snitch_regfile.mem[218] ),
    .A3(\i_snitch.i_snitch_regfile.mem[250] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1  (.S0(net2999),
    .A0(\i_snitch.i_snitch_regfile.mem[154] ),
    .A1(\i_snitch.i_snitch_regfile.mem[186] ),
    .A2(\i_snitch.i_snitch_regfile.mem[218] ),
    .A3(\i_snitch.i_snitch_regfile.mem[250] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[122]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net3085),
    .C1(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2849),
    .A1(net3075),
    .Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2751));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net887),
    .A2(net2445),
    .A1(net2252));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3192),
    .D(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[155] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2885),
    .B(net2657));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[155] ),
    .A1(\i_snitch.i_snitch_regfile.mem[187] ),
    .A2(\i_snitch.i_snitch_regfile.mem[219] ),
    .A3(\i_snitch.i_snitch_regfile.mem[251] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1  (.S0(net2999),
    .A0(\i_snitch.i_snitch_regfile.mem[155] ),
    .A1(\i_snitch.i_snitch_regfile.mem[187] ),
    .A2(\i_snitch.i_snitch_regfile.mem[219] ),
    .A3(\i_snitch.i_snitch_regfile.mem[251] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[123]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2836),
    .A2(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net3084),
    .C1(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2849),
    .A1(net3075),
    .Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2751));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2816),
    .B(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2349),
    .B2(net937),
    .A2(net2447),
    .A1(net2246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[156] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2886),
    .B(net2655));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0  (.S0(net3119),
    .A0(\i_snitch.i_snitch_regfile.mem[156] ),
    .A1(\i_snitch.i_snitch_regfile.mem[188] ),
    .A2(\i_snitch.i_snitch_regfile.mem[220] ),
    .A3(\i_snitch.i_snitch_regfile.mem[252] ),
    .S1(net3100),
    .X(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1  (.S0(net3004),
    .A0(\i_snitch.i_snitch_regfile.mem[156] ),
    .A1(\i_snitch.i_snitch_regfile.mem[188] ),
    .A2(\i_snitch.i_snitch_regfile.mem[220] ),
    .A3(\i_snitch.i_snitch_regfile.mem[252] ),
    .S1(net2978),
    .X(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2837),
    .A2(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2817),
    .A2(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net1098),
    .A2(net2446),
    .A1(net2250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[157] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2889),
    .B(net2653));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0  (.S0(net3126),
    .A0(\i_snitch.i_snitch_regfile.mem[157] ),
    .A1(\i_snitch.i_snitch_regfile.mem[189] ),
    .A2(\i_snitch.i_snitch_regfile.mem[221] ),
    .A3(\i_snitch.i_snitch_regfile.mem[253] ),
    .S1(net3106),
    .X(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1  (.S0(net3012),
    .A0(\i_snitch.i_snitch_regfile.mem[157] ),
    .A1(\i_snitch.i_snitch_regfile.mem[189] ),
    .A2(\i_snitch.i_snitch_regfile.mem[221] ),
    .A3(\i_snitch.i_snitch_regfile.mem[253] ),
    .S1(net2985),
    .X(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[125]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2639),
    .B(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net3080),
    .C1(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(net2850),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2753));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2351),
    .B2(net971),
    .A2(net2446),
    .A1(net2244));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[158] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2889),
    .B(net2649));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0  (.S0(net3126),
    .A0(\i_snitch.i_snitch_regfile.mem[158] ),
    .A1(\i_snitch.i_snitch_regfile.mem[190] ),
    .A2(\i_snitch.i_snitch_regfile.mem[222] ),
    .A3(\i_snitch.i_snitch_regfile.mem[254] ),
    .S1(net3106),
    .X(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1  (.S0(net3012),
    .A0(\i_snitch.i_snitch_regfile.mem[158] ),
    .A1(\i_snitch.i_snitch_regfile.mem[190] ),
    .A2(\i_snitch.i_snitch_regfile.mem[222] ),
    .A3(\i_snitch.i_snitch_regfile.mem[254] ),
    .S1(net2985),
    .X(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2838),
    .A2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B  (.A(net2639),
    .B(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1  (.A1(net3078),
    .A2(net2850),
    .Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_A ),
    .A(net3074),
    .B(net2753));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B  (.A(net2819),
    .B(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2349),
    .B2(net924),
    .A2(net2645),
    .A1(net2887));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[159] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2347));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0  (.S0(net3124),
    .A0(\i_snitch.i_snitch_regfile.mem[159] ),
    .A1(\i_snitch.i_snitch_regfile.mem[191] ),
    .A2(\i_snitch.i_snitch_regfile.mem[223] ),
    .A3(\i_snitch.i_snitch_regfile.mem[255] ),
    .S1(net3103),
    .X(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1  (.S0(net3009),
    .A0(\i_snitch.i_snitch_regfile.mem[159] ),
    .A1(\i_snitch.i_snitch_regfile.mem[191] ),
    .A2(\i_snitch.i_snitch_regfile.mem[223] ),
    .A3(\i_snitch.i_snitch_regfile.mem[255] ),
    .S1(net2982),
    .X(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[127]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2837),
    .A2(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C  (.A(net2642),
    .B(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1  (.A2(net2720),
    .A1(net3074),
    .B1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B  (.A(net2701),
    .B(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2818),
    .A2(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[160]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2343),
    .B2(net910),
    .A2(net2903),
    .A1(net2773));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[160] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[160]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2340));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[161] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2443),
    .B2(net2514),
    .A2(net2902),
    .A1(net2773));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[161]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net464),
    .B(net2342));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[161]_sg13g2_nand2_1_A_1  (.Y(\i_snitch.i_snitch_regfile.mem[161]_sg13g2_nand2_1_A_1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[161] ),
    .B(net2826));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[162] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2442),
    .A1(net2771),
    .Y(\i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[162]_sg13g2_nor3_1_A  (.A(net1282),
    .B(net2772),
    .C(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[162]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[163] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2443),
    .A1(net2772),
    .Y(\i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[163]_sg13g2_nor3_1_A  (.A(net1309),
    .B(net2772),
    .C(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[163]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[164] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2442),
    .A1(net2773),
    .Y(\i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[164]_sg13g2_nor3_1_A  (.A(net1290),
    .B(net2776),
    .C(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[164]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[165] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2442),
    .A1(net2771),
    .Y(\i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[165]_sg13g2_nor3_1_A  (.A(net1239),
    .B(net2772),
    .C(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[165]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[166]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2344),
    .B2(net1135),
    .A2(net2899),
    .A1(net2774));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[166] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[166]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2444));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[167]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2442),
    .B2(net2284),
    .A2(net2342),
    .A1(net1163));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[167] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[167]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2771),
    .B(net2897));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[168]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2343),
    .B2(net953),
    .A2(net2643),
    .A1(net2773));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[168] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[168]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[169]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2343),
    .B2(net1029),
    .A2(net2686),
    .A1(net2773));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[169] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[169]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[170]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .B2(net2282),
    .A2(net2344),
    .A1(net1192));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3278),
    .D(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[170] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[170]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2774),
    .B(net2693));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[171]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net897),
    .A2(net2679),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[171] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[171]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[172]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net705),
    .A2(net2692),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[172] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[172]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[173]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2344),
    .B2(net1002),
    .A2(net2690),
    .A1(net2774));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[173] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[173]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2444));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[174]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2344),
    .B2(net974),
    .A2(net2688),
    .A1(net2774));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[174] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[174]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2444));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[175]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net906),
    .A2(net2678),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[175] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[175]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[176]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2444),
    .B2(net2263),
    .A2(net2344),
    .A1(net1275));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[176] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[176]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2774),
    .B(net2668));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[177]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net727),
    .A2(net2664),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[177] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[177]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[178]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2444),
    .B2(net2272),
    .A2(net2344),
    .A1(net1178));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[178] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[178]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2774),
    .B(net2675));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[179]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2442),
    .B2(net2270),
    .A2(net2342),
    .A1(net1259));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[179] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[179]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2771),
    .B(net2673));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[180]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net866),
    .A2(net2671),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[180] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[180]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2341));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[181]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2443),
    .B2(net2268),
    .A2(net2342),
    .A1(net1175));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[181] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[181]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2772),
    .B(net2669));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[182]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net1045),
    .A2(net2651),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[182] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[182]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2341));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[183]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net1078),
    .A2(net2648),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[183] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[183]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2341));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[184]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2345),
    .B2(net790),
    .A2(net2665),
    .A1(net2775));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[184] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[184]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2341));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[185]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2442),
    .B2(net2266),
    .A2(net2342),
    .A1(net1188));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[185] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[185]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2771),
    .B(net2661));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[186]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2442),
    .B2(net2254),
    .A2(net2342),
    .A1(net1215));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[186] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[186]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2771),
    .B(net2659));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[187]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2442),
    .B2(net2252),
    .A2(net2342),
    .A1(net1278));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3192),
    .D(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[187] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[187]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2771),
    .B(net2657));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[188]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2443),
    .B2(net2246),
    .A2(net2342),
    .A1(net1190));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[188] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[188]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2772),
    .B(net2655));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[189]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2444),
    .B2(net2250),
    .A2(net2344),
    .A1(net1276));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[189] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[189]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2774),
    .B(net2653));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[190]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .B2(net2244),
    .A2(net2344),
    .A1(net1244));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[190] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[190]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2774),
    .B(net2649));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[191]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2343),
    .B2(net840),
    .A2(net2645),
    .A1(net2773));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[191] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[191]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2340));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[192]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2339),
    .B2(net1048),
    .A2(net2903),
    .A1(net2790));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[192] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[192]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2334));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[193] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2440),
    .B2(net2513),
    .A2(net2901),
    .A1(net2791));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[193] ),
    .A1(\i_snitch.i_snitch_regfile.mem[225] ),
    .S(net3013),
    .X(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_X ));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_1  (.A0(\i_snitch.i_snitch_regfile.mem[193] ),
    .A1(\i_snitch.i_snitch_regfile.mem[225] ),
    .S(net3133),
    .X(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_1_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[193]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net452),
    .B(net2337));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[194] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2439),
    .A1(net2788),
    .Y(\i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[194]_sg13g2_nor3_1_A  (.A(net1238),
    .B(net2788),
    .C(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[194]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[195] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2441),
    .A1(net2789),
    .Y(\i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[195]_sg13g2_nor3_1_A  (.A(net1360),
    .B(net2789),
    .C(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[195]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[196] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2439),
    .A1(net2790),
    .Y(\i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[196]_sg13g2_nor3_1_A  (.A(net1329),
    .B(net2790),
    .C(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[196]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[197] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2439),
    .A1(net2788),
    .Y(\i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[197]_sg13g2_nor3_1_A  (.A(net1312),
    .B(net2789),
    .C(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[197]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[198]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2337),
    .B2(net1113),
    .A2(net2900),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[198] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[198]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2440));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[199]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net885),
    .A2(net2439),
    .A1(net2284));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[199] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[199]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2788),
    .B(net2897));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[200]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net823),
    .A2(net2643),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[200] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[200]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[201]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2339),
    .B2(net739),
    .A2(net2686),
    .A1(net2790));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[201] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[201]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[202]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net913),
    .A2(net2440),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3278),
    .D(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[202] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[202]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2792),
    .B(net2693));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[203]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2339),
    .B2(net870),
    .A2(net2679),
    .A1(net2793));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[203] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[203]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[204]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net926),
    .A2(net2692),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[204] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[204]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[205]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net1041),
    .A2(net2690),
    .A1(net2792));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[205] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[205]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2440));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[206]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net1084),
    .A2(net2688),
    .A1(net2792));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3289),
    .D(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[206] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[206]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2440));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[207]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2339),
    .B2(net1080),
    .A2(net2678),
    .A1(net2793));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[207] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[207]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[208]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net980),
    .A2(net2441),
    .A1(net2263));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3289),
    .D(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[208] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[208]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2792),
    .B(net2668));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[209]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2339),
    .B2(net1039),
    .A2(net2664),
    .A1(net2793));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[209] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[209]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[210]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net968),
    .A2(net2441),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[210] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[210]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2792),
    .B(net2675));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[211]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net863),
    .A2(net2439),
    .A1(net2270));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[211] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[211]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2788),
    .B(net2673));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[212]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net718),
    .A2(net2671),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3323),
    .D(\i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[212] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[212]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2335));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[213]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net1132),
    .A2(net2441),
    .A1(net2268));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[213] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[213]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2789),
    .B(net2669));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[214]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net1106),
    .A2(net2651),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[214] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[214]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2335));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[215]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net791),
    .A2(net2648),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[215] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[215]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2335));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[216]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2337),
    .B2(net808),
    .A2(net2666),
    .A1(net2791));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[216] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[216]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2335),
    .A2(net2257));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[217]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net857),
    .A2(net2439),
    .A1(net2266));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[217] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[217]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2788),
    .B(net2661));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[218]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net1092),
    .A2(net2439),
    .A1(net2254));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[218] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[218]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2788),
    .B(net2659));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[219]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net984),
    .A2(net2439),
    .A1(net2252));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[219] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[219]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2788),
    .B(net2657));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[220]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2336),
    .B2(net970),
    .A2(net2440),
    .A1(net2246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[220] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[220]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2789),
    .B(net2655));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[221]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net1016),
    .A2(net2440),
    .A1(net2250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[221] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[221]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2792),
    .B(net2653));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[222]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2338),
    .B2(net972),
    .A2(net2440),
    .A1(net2244));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3271),
    .D(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[222] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[222]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2792),
    .B(net2649));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[223]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2336),
    .B2(net756),
    .A2(net2646),
    .A1(net2790));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3305),
    .D(\i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[223] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[223]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2334));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[224]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2333),
    .B2(net783),
    .A2(net2903),
    .A1(net2874));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[224] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[224]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2328));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[225] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2437),
    .B2(net2513),
    .A2(net2901),
    .A1(net2875));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[225]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[225]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net444),
    .B(net2331));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[226] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2436),
    .A1(net2872),
    .Y(\i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[226]_sg13g2_nor3_1_A  (.A(net1357),
    .B(net2872),
    .C(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[226]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[227] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2478),
    .C1(\i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2436),
    .A1(net2873),
    .Y(\i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[227]_sg13g2_nor3_1_A  (.A(net1327),
    .B(net2873),
    .C(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[227]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[228] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2436),
    .A1(net2874),
    .Y(\i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[228]_sg13g2_nor3_1_A  (.A(net1338),
    .B(net2874),
    .C(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[228]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[229] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2436),
    .A1(net2872),
    .Y(\i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[229]_sg13g2_nor3_1_A  (.A(net1368),
    .B(net2872),
    .C(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[229]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[230]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net918),
    .A2(net2900),
    .A1(net2876));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[230] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[230]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2437));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[231]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net1064),
    .A2(net2436),
    .A1(net2284));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[231] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[231]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2873),
    .B(net2897));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[232]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net1137),
    .A2(net2643),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[232] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[232]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[233]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2333),
    .B2(net1032),
    .A2(net2686),
    .A1(net2874));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[233] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[233]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[234]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net1028),
    .A2(net2437),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3278),
    .D(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[234] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[234]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2876),
    .B(net2693));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[235]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net896),
    .A2(net2679),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[235] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[235]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[236]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net1056),
    .A2(net2692),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[236] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[236]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[237]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net1144),
    .A2(net2690),
    .A1(net2876));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[237] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[237]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2437));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[238]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net835),
    .A2(net2688),
    .A1(net2876));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[238] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[238]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2437));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[239]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2333),
    .B2(net1128),
    .A2(net2677),
    .A1(net2877));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3299),
    .D(\i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[239] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[239]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[240]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net1058),
    .A2(net2438),
    .A1(net2263));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3289),
    .D(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[240] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[240]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2876),
    .B(net2668));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[241]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2333),
    .B2(net979),
    .A2(net2664),
    .A1(net2877));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[241] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[241]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[242]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net1012),
    .A2(net2438),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[242] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[242]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2876),
    .B(net2675));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[243]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net1023),
    .A2(net2436),
    .A1(net2270));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[243] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[243]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2872),
    .B(net2673));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[244]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net724),
    .A2(net2671),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3323),
    .D(\i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[244] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[244]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2329));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[245]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net1095),
    .A2(net2438),
    .A1(net2268));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[245] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[245]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2873),
    .B(net2669));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[246]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net903),
    .A2(net2651),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3320),
    .D(\i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[246] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[246]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2329));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[247]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net1005),
    .A2(net2648),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[247] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[247]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2329));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[248]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2331),
    .B2(net899),
    .A2(net2666),
    .A1(net2875));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[248] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[248]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2329),
    .A2(net2257));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[249]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net1006),
    .A2(net2438),
    .A1(net2266));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[249] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[249]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2872),
    .B(net2661));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[250]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net993),
    .A2(net2436),
    .A1(net2254));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3207),
    .D(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[250] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[250]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2872),
    .B(net2659));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[251]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net782),
    .A2(net2436),
    .A1(net2252));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[251] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[251]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2872),
    .B(net2657));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[252]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2330),
    .B2(net1024),
    .A2(net2437),
    .A1(net2246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[252] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[252]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2873),
    .B(net2655));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[253]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net958),
    .A2(net2437),
    .A1(net2250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3271),
    .D(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[253] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[253]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2876),
    .B(net2653));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[254]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2332),
    .B2(net921),
    .A2(net2437),
    .A1(net2244));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[254] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[254]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2876),
    .B(net2649));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[255]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2330),
    .B2(net761),
    .A2(net2646),
    .A1(net2874));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3305),
    .D(\i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[255] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[255]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2328));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2323),
    .B2(net865),
    .A2(net2904),
    .A1(net2892));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3255),
    .D(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[256] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2322));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[256] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2919));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(net2931),
    .B(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0  (.S0(net3010),
    .A0(\i_snitch.i_snitch_regfile.mem[256] ),
    .A1(\i_snitch.i_snitch_regfile.mem[288] ),
    .A2(\i_snitch.i_snitch_regfile.mem[320] ),
    .A3(\i_snitch.i_snitch_regfile.mem[352] ),
    .S1(net2983),
    .X(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ),
    .C1(net2957),
    .B1(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2969),
    .Y(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[257] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2434),
    .B2(net2514),
    .A2(net2902),
    .A1(net2894));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0  (.S0(net3013),
    .A0(\i_snitch.i_snitch_regfile.mem[257] ),
    .A1(\i_snitch.i_snitch_regfile.mem[289] ),
    .A2(\i_snitch.i_snitch_regfile.mem[385] ),
    .A3(\i_snitch.i_snitch_regfile.mem[417] ),
    .S1(net2963),
    .X(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2954),
    .A2(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C  (.A(net2640),
    .B(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1  (.B2(net2981),
    .C1(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ),
    .A1(net3104),
    .Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2752));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[257]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net505),
    .B(net2324));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[258] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net701),
    .C1(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2327),
    .A1(net2485),
    .Y(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2435));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2891),
    .B(net2912),
    .X(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[258] ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[259] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2478),
    .C1(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2433),
    .A1(net2892),
    .Y(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[259]_sg13g2_nor3_1_A  (.A(net1359),
    .B(net2892),
    .C(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[259] ),
    .A2(net2814));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ),
    .A(net2942),
    .B(net2953));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[260] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net693),
    .C1(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2327),
    .A1(net2892),
    .Y(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2476),
    .B(net2433),
    .X(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[260] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y ),
    .A2(net3007));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0  (.S0(net3122),
    .A0(\i_snitch.i_snitch_regfile.mem[260] ),
    .A1(\i_snitch.i_snitch_regfile.mem[292] ),
    .A2(\i_snitch.i_snitch_regfile.mem[324] ),
    .A3(\i_snitch.i_snitch_regfile.mem[356] ),
    .S1(net3104),
    .X(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X ),
    .A1(net2939),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[261] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net673),
    .C1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2323),
    .A1(net2408),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2435));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2891),
    .B(net2906),
    .X(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[261] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y ),
    .A2(net3001));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0  (.S0(net3118),
    .A0(\i_snitch.i_snitch_regfile.mem[261] ),
    .A1(\i_snitch.i_snitch_regfile.mem[293] ),
    .A2(\i_snitch.i_snitch_regfile.mem[325] ),
    .A3(\i_snitch.i_snitch_regfile.mem[357] ),
    .S1(net3102),
    .X(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2935),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A1(net3089),
    .B1(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B  (.A(net2634),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2b_2 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y_sg13g2_nor2b_1_A  (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_B_Y ),
    .B_N(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ),
    .B2(net3087),
    .A2(net2719),
    .A1(\i_req_arb.data_i[40] ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B  (.A(net2579),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2  (.A1(net60),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(net2564));
 sg13g2_and4_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D  (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .B(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ),
    .D(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X ));
 sg13g2_nor4_2 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A_sg13g2_nor4_1_Y  (.A(net2608),
    .B(net2593),
    .C(net2561),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .D(net2589));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X ),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y ),
    .B1(net2565));
 sg13g2_xnor2_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y_sg13g2_xnor2_1_B  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_a21oi_1_A1_Y ));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B  (.B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X ),
    .C(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C ),
    .A(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C_sg13g2_inv_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_B_C ),
    .A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X_sg13g2_nor2_1_B  (.A(net2565),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_X ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D  (.B(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor4_2 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D  (.A(net2579),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B ),
    .C(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B_sg13g2_a21oi_1_A2  (.A1(net2570),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .B1(net2579));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B_sg13g2_nand4_1_Y  (.B(net2599),
    .C(net2556),
    .A(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B ),
    .D(net2602));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2  (.B1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2564),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y ));
 sg13g2_or3_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C  (.A(net2564),
    .B(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2325),
    .B2(net1150),
    .A2(net2899),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[262] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2435));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[262] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2920));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0  (.S0(net3014),
    .A0(\i_snitch.i_snitch_regfile.mem[262] ),
    .A1(\i_snitch.i_snitch_regfile.mem[294] ),
    .A2(\i_snitch.i_snitch_regfile.mem[326] ),
    .A3(\i_snitch.i_snitch_regfile.mem[358] ),
    .S1(net2986),
    .X(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2958),
    .B1(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2639),
    .B(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1  (.A2(net2752),
    .A1(net3086),
    .B1(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2323),
    .B2(net1114),
    .A2(net2433),
    .A1(net2284));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[263] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2898));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[263] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y ),
    .A2(net3002));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_mux4_1_A0  (.S0(net3118),
    .A0(\i_snitch.i_snitch_regfile.mem[263] ),
    .A1(\i_snitch.i_snitch_regfile.mem[295] ),
    .A2(\i_snitch.i_snitch_regfile.mem[327] ),
    .A3(\i_snitch.i_snitch_regfile.mem[359] ),
    .S1(net3099),
    .X(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[263]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2935),
    .A2(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_mux4_1_A0_X ),
    .Y(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2325),
    .B2(net634),
    .A2(net2644),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3308),
    .D(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[264] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2321));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[264] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y ),
    .A2(net110),
    .Y(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y ),
    .A2(net3019));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2327),
    .B2(net644),
    .A2(net2685),
    .A1(net2892));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[265] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2322));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[265] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2919));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1  (.A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1  (.B2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ),
    .C1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(net3080),
    .A1(\i_req_arb.data_i[44] ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2720));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y ),
    .A2(net3008));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net1020),
    .A2(net2434),
    .A1(net2283));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[266] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2694));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[266] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2920));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0  (.S0(net3013),
    .A0(\i_snitch.i_snitch_regfile.mem[266] ),
    .A1(\i_snitch.i_snitch_regfile.mem[298] ),
    .A2(\i_snitch.i_snitch_regfile.mem[330] ),
    .A3(\i_snitch.i_snitch_regfile.mem[362] ),
    .S1(net2986),
    .X(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2970),
    .A2(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2325),
    .B2(net787),
    .A2(net2680),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[267] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2321));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[267] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y ),
    .A2(net3020));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0  (.S0(net3135),
    .A0(\i_snitch.i_snitch_regfile.mem[267] ),
    .A1(\i_snitch.i_snitch_regfile.mem[299] ),
    .A2(\i_snitch.i_snitch_regfile.mem[331] ),
    .A3(\i_snitch.i_snitch_regfile.mem[363] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X ),
    .A1(net2937),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[268]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[268] ),
    .A2(net3029),
    .Y(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2991));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[268]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2326),
    .B2(net811),
    .A2(net2691),
    .A1(net2894));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3308),
    .D(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[268] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2321));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[268]_sg13g2_o21ai_1_A1  (.B1(net2937),
    .Y(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[268] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2324),
    .B2(net704),
    .A2(net2689),
    .A1(net2895));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[269] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2434));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[269] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2920));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2632),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2724),
    .A1(\i_snitch.inst_addr_o[13] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y ),
    .A2(net3017));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[270] ),
    .A2(net3028),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2988));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net940),
    .A2(net2687),
    .A1(net2895));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[270] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2435));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[270] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2920));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2631),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2725),
    .A1(\i_snitch.inst_addr_o[14] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[271]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[271] ),
    .A2(net3029),
    .Y(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[271]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2326),
    .B2(net1030),
    .A2(net2677),
    .A1(net2894));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[271] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2321));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[271]_sg13g2_o21ai_1_A1  (.B1(net2937),
    .Y(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[271] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net1229),
    .A2(net2434),
    .A1(net2263));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[272] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2668));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[272] ),
    .B(net3028));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[272]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[272] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2325),
    .B2(net562),
    .A2(net2663),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[273] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2321));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[273] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2920));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y ),
    .C1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ),
    .B1(net2637),
    .A1(\i_snitch.inst_addr_o[17] ),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net2724));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y ),
    .A2(net3020));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[274] ),
    .A2(net3028),
    .Y(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2987));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net989),
    .A2(net2434),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3287),
    .D(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[274] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2676));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[274]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[274] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2323),
    .B2(net1143),
    .A2(net2433),
    .A1(net2270));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[275] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2673));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[275] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2918));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0  (.S0(net3000),
    .A0(\i_snitch.i_snitch_regfile.mem[275] ),
    .A1(\i_snitch.i_snitch_regfile.mem[307] ),
    .A2(\i_snitch.i_snitch_regfile.mem[339] ),
    .A3(\i_snitch.i_snitch_regfile.mem[371] ),
    .S1(net2976),
    .X(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2968),
    .A2(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[276]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[276] ),
    .A2(net3030),
    .Y(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2993));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[276]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2325),
    .B2(net785),
    .A2(net2672),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3315),
    .D(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[276] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2321));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[276]_sg13g2_o21ai_1_A1  (.B1(net2937),
    .Y(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[276] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2323),
    .B2(net691),
    .A2(net2433),
    .A1(net2269));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3264),
    .D(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[277] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2670));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[277] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y ),
    .A2(net2918),
    .Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net3092));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y ),
    .A2(net3005));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2325),
    .B2(net944),
    .A2(net2652),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[278] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2321));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0  (.S0(net3133),
    .A0(\i_snitch.i_snitch_regfile.mem[278] ),
    .A1(\i_snitch.i_snitch_regfile.mem[310] ),
    .A2(\i_snitch.i_snitch_regfile.mem[342] ),
    .A3(\i_snitch.i_snitch_regfile.mem[374] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X ),
    .A1(net2938),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[278]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[278] ),
    .B(net3029));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2325),
    .B2(net912),
    .A2(net2647),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[279] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2321));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[279] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y ),
    .A2(net3019));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0  (.S0(net3134),
    .A0(\i_snitch.i_snitch_regfile.mem[279] ),
    .A1(\i_snitch.i_snitch_regfile.mem[311] ),
    .A2(\i_snitch.i_snitch_regfile.mem[343] ),
    .A3(\i_snitch.i_snitch_regfile.mem[375] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X ),
    .A1(net2938),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[280]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2325),
    .B2(net1118),
    .A2(net2666),
    .A1(net2893));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3315),
    .D(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[280] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net310),
    .A2(net2322));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[280]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[280] ),
    .B(net3029));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[280]_sg13g2_o21ai_1_A1  (.B1(net2938),
    .Y(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[280] ),
    .A2(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2323),
    .B2(net700),
    .A2(net2433),
    .A1(net2267));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3216),
    .D(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[281] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2662));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[281] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2918));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2721),
    .A1(\i_snitch.inst_addr_o[25] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y ),
    .A2(net3004));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2323),
    .B2(net683),
    .A2(net2433),
    .A1(net2254));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3208),
    .D(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[282] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2660));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[282] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y ),
    .A2(net2918),
    .Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y ),
    .A2(net3000));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2323),
    .B2(net670),
    .A2(net2433),
    .A1(net2252));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[283] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2891),
    .B(net2657));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[283] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(net3098),
    .C1(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2918));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2509),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2720),
    .A1(\i_snitch.inst_addr_o[27] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y ),
    .A2(net2999));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net1067),
    .A2(net2434),
    .A1(net2247));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[284] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2655));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0  (.S0(net3005),
    .A0(\i_snitch.i_snitch_regfile.mem[284] ),
    .A1(\i_snitch.i_snitch_regfile.mem[316] ),
    .A2(\i_snitch.i_snitch_regfile.mem[348] ),
    .A3(\i_snitch.i_snitch_regfile.mem[380] ),
    .S1(net2977),
    .X(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2958),
    .B1(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1  (.B2(net3082),
    .C1(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .B1(net2850),
    .A1(net3074),
    .Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2754));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[284]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[284] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2324),
    .B2(net884),
    .A2(net2434),
    .A1(net2251));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[285] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2654));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0  (.S0(net3126),
    .A0(\i_snitch.i_snitch_regfile.mem[285] ),
    .A1(\i_snitch.i_snitch_regfile.mem[317] ),
    .A2(\i_snitch.i_snitch_regfile.mem[349] ),
    .A3(\i_snitch.i_snitch_regfile.mem[381] ),
    .S1(net3106),
    .X(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X ),
    .A1(net2936),
    .B1(net2930),
    .X(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[285]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[285] ),
    .B(net3028));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2327),
    .B2(net671),
    .A2(net2434),
    .A1(net2245));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[286] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2895),
    .B(net2650));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[286] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2921));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.inst_addr_o[30] ),
    .A2(net2721),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_B1 ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y ),
    .A2(net3012));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2326),
    .B2(net917),
    .A2(net2645),
    .A1(net2894));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[287] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2322));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0  (.S0(net3123),
    .A0(\i_snitch.i_snitch_regfile.mem[287] ),
    .A1(\i_snitch.i_snitch_regfile.mem[319] ),
    .A2(\i_snitch.i_snitch_regfile.mem[351] ),
    .A3(\i_snitch.i_snitch_regfile.mem[383] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1  (.S0(net3008),
    .A0(\i_snitch.i_snitch_regfile.mem[287] ),
    .A1(\i_snitch.i_snitch_regfile.mem[319] ),
    .A2(\i_snitch.i_snitch_regfile.mem[351] ),
    .A3(\i_snitch.i_snitch_regfile.mem[383] ),
    .S1(net2982),
    .X(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ),
    .C1(net2957),
    .B1(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2969),
    .Y(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net2937),
    .A2(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(net2932));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[288]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2904),
    .B2(net2778),
    .A2(net2316),
    .A1(net1254));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3255),
    .D(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[288] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2315),
    .A2(net2522));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[288]_sg13g2_o21ai_1_A1  (.B1(net2939),
    .Y(\i_snitch.i_snitch_regfile.mem[288]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[288] ),
    .A2(net2811));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[289]_sg13g2_a221oi_1_A1  (.B2(net2920),
    .C1(net3094),
    .B1(\i_snitch.i_snitch_regfile.mem[257] ),
    .A1(\i_snitch.i_snitch_regfile.mem[289] ),
    .Y(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2825));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[289]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2901),
    .B2(net2779),
    .A2(net2317),
    .A1(net1316));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[289] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2431),
    .B(net2513));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[290] ),
    .A2(net3002),
    .Y(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2975));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A_Y ),
    .A2(net3002));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[290] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2485),
    .C1(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2430),
    .A1(net657),
    .Y(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2316));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2777),
    .B(net2912),
    .X(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[290] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A_Y ),
    .C1(net3091),
    .B1(net2918),
    .A1(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2825));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[291] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2778),
    .C1(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2910),
    .A1(net678),
    .Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2320));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2432),
    .B(net2478),
    .X(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[291] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2825));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1  (.S0(net3006),
    .A0(\i_snitch.i_snitch_regfile.mem[259] ),
    .A1(\i_snitch.i_snitch_regfile.mem[291] ),
    .A2(\i_snitch.i_snitch_regfile.mem[323] ),
    .A3(\i_snitch.i_snitch_regfile.mem[355] ),
    .S1(net2979),
    .X(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2640),
    .B(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2b_2 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ),
    .B2(net2955),
    .A2(net2752),
    .A1(net3089));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[292]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[292] ),
    .A2(net3007),
    .Y(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2980));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[292] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2778),
    .C1(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2908),
    .A1(net2430),
    .Y(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2476));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[292]_sg13g2_nor3_1_A  (.A(net1320),
    .B(net2778),
    .C(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[292]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[293]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[293] ),
    .A2(net3001),
    .Y(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2975));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[293] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2777),
    .C1(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2906),
    .A1(net2430),
    .Y(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2408));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[293]_sg13g2_nor3_1_A  (.A(net1304),
    .B(net2777),
    .C(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[293]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[294]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2899),
    .B2(net2779),
    .A2(net2317),
    .A1(net1209));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[294] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2431),
    .B(net2287));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[294]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[294]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[294] ),
    .A2(net2812));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[295]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[295] ),
    .A2(net3002),
    .Y(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2975));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[295]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2430),
    .B2(net2285),
    .A2(net2316),
    .A1(net1218));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[295] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[295]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2777),
    .B(net2898));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[296]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[296] ),
    .A2(net3019),
    .Y(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[296]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2643),
    .B2(net2780),
    .A2(net2318),
    .A1(net1318));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3308),
    .D(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[296] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2279));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[296]_sg13g2_o21ai_1_A1  (.B1(net2937),
    .Y(\i_snitch.i_snitch_regfile.mem[296]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[296] ),
    .A2(net2813));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[297]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[297] ),
    .A2(net3008),
    .Y(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2982));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[297]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2685),
    .B2(net2778),
    .A2(net2320),
    .A1(net1280));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[297] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2315),
    .A2(net2299));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[297]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[297]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[297] ),
    .A2(net2811));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[298]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2431),
    .B2(net2283),
    .A2(net2317),
    .A1(net1257));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[298] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2779),
    .B(net2694));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[298]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[298]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[298] ),
    .A2(net2812));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[299]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[299] ),
    .A2(net3021),
    .Y(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[299]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2680),
    .B2(net2780),
    .A2(net2318),
    .A1(net1351));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[299] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[299]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2281));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2691),
    .B2(net2780),
    .A2(net2318),
    .A1(net1138));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[300] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2276));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[300] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2829));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2632),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2724),
    .A1(\i_snitch.inst_addr_o[12] ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[300]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[300] ),
    .B(net3024));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[301] ),
    .A2(net3017),
    .Y(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2988));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2689),
    .B2(net2779),
    .A2(net2317),
    .A1(net1260));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[301] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2431),
    .B(net2291));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[301]_sg13g2_o21ai_1_A1  (.B1(net2938),
    .Y(\i_snitch.i_snitch_regfile.mem[301]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[301] ),
    .A2(net2812));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2687),
    .B2(net2779),
    .A2(net2317),
    .A1(net1231));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[302] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2431),
    .B(net2275));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[302] ),
    .B(net3017));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[302]_sg13g2_o21ai_1_A1  (.B1(net2938),
    .Y(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[302] ),
    .A2(net2812));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2677),
    .B2(net2781),
    .A2(net2319),
    .A1(net1081));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[303] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2264));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[303] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y ),
    .A2(net2829),
    .Y(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[271]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y ),
    .A2(net3029));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[304] ),
    .A2(net3016),
    .Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2987));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2431),
    .B2(net2263),
    .A2(net2317),
    .A1(net1243));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3286),
    .D(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[304] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2779),
    .B(net2668));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[304] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_nand2_1_A_1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2827));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2511),
    .Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2632),
    .Y(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1  (.A2(net2725),
    .A1(\i_snitch.inst_addr_o[16] ),
    .B1(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[305]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[305] ),
    .A2(net3020),
    .Y(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2992));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[305]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2663),
    .B2(net2781),
    .A2(net2319),
    .A1(net1266));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[305] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2288));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[305]_sg13g2_o21ai_1_A1  (.B1(net2937),
    .Y(\i_snitch.i_snitch_regfile.mem[305]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[305] ),
    .A2(net2812));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[306] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2676),
    .B2(net2781),
    .A2(net2273),
    .A1(net2432));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[306] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y ),
    .A2(net2827),
    .Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net456),
    .B(net2319));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[306]_sg13g2_nand2_1_A_1  (.Y(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_nand2_1_A_1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[306] ),
    .B(net3016));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[307]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2430),
    .B2(net2271),
    .A2(net2316),
    .A1(net1292));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[307] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2777),
    .B(net2674));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[307]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[307]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[307] ),
    .A2(net2810));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2672),
    .B2(net2780),
    .A2(net2318),
    .A1(net1195));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3316),
    .D(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[308] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2261));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[308] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2828));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2632),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2636),
    .A2(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2722),
    .A1(\i_snitch.inst_addr_o[20] ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[308]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[308] ),
    .B(net3020));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[309] ),
    .A2(net3005),
    .Y(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2978));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2432),
    .B2(net2269),
    .A2(net2316),
    .A1(net1221));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[309] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2778),
    .B(net2670));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[309]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[309] ),
    .A2(net2810));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[310]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[310] ),
    .A2(net3020),
    .Y(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[310]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2652),
    .B2(net2780),
    .A2(net2318),
    .A1(net1152));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[310] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2259));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[311]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[311] ),
    .A2(net3019),
    .Y(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2991));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[311]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2647),
    .B2(net2780),
    .A2(net2318),
    .A1(net1182));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3310),
    .D(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[311] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[311]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2314),
    .A2(net2248));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[312] ),
    .A2(net3022),
    .Y(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2666),
    .B2(net2780),
    .A2(net2318),
    .A1(net1246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[312] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2315),
    .A2(net310));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[312] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y ),
    .A2(net2828),
    .Y(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[313] ),
    .A2(net3004),
    .Y(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2977));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2430),
    .B2(net2267),
    .A2(net2316),
    .A1(net1268));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[313] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2777),
    .B(net2662));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[313]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[313]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[313] ),
    .A2(net2810));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[314] ),
    .A2(net3000),
    .Y(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2976));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2430),
    .B2(net2255),
    .A2(net2316),
    .A1(net1205));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3208),
    .D(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[314] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2777),
    .B(net2660));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[314]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[314]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[314] ),
    .A2(net2810));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[315] ),
    .A2(net2999),
    .Y(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2973));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2430),
    .B2(net2253),
    .A2(net2316),
    .A1(net1162));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[315] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2777),
    .B(net2658));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[315]_sg13g2_o21ai_1_A1  (.B1(net2935),
    .Y(\i_snitch.i_snitch_regfile.mem[315]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[315] ),
    .A2(net2810));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2431),
    .B2(net2247),
    .A2(net2317),
    .A1(net1171));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[316] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2779),
    .B(net2656));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[316] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2825));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[317]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[317] ),
    .A2(net3012),
    .Y(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2985));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[317]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2431),
    .B2(net2251),
    .A2(net2317),
    .A1(net1211));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[317] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2779),
    .B(net2654));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[318] ),
    .A2(net3015),
    .Y(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2986));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2432),
    .B2(net2245),
    .A2(net2319),
    .A1(net1161));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[318] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2781),
    .B(net2650));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[318]_sg13g2_o21ai_1_A1  (.B1(net2936),
    .Y(\i_snitch.i_snitch_regfile.mem[318]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[318] ),
    .A2(net2812));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[319]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2645),
    .B2(net2780),
    .A2(net2318),
    .A1(net1232));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[319] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[319]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2315),
    .A2(net2242));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[320]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2402),
    .B2(net717),
    .A2(net2904),
    .A1(net2795));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3255),
    .D(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[320] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2400));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[320]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[320]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[320] ),
    .B(net2949));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[321] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2473),
    .B2(net2513),
    .A2(net2901),
    .A1(net2796));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0  (.S0(net3013),
    .A0(\i_snitch.i_snitch_regfile.mem[321] ),
    .A1(\i_snitch.i_snitch_regfile.mem[353] ),
    .A2(\i_snitch.i_snitch_regfile.mem[449] ),
    .A3(\i_snitch.i_snitch_regfile.mem[481] ),
    .S1(net2963),
    .X(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .C1(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[193]_sg13g2_mux2_1_A0_X ),
    .A1(net2954),
    .Y(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_mux4_1_A0_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net470),
    .B(net2403));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_o21ai_1_A1  (.B1(net3107),
    .Y(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[321] ),
    .A2(net3128));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[321]_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_B1 ),
    .A(\i_snitch.i_snitch_regfile.mem[321]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[322] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net690),
    .C1(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2402),
    .A1(net2485),
    .Y(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2474));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2795),
    .B(net2912),
    .X(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[322] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[322] ),
    .B(net2947));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B  (.B(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_nand2_1_A_Y ),
    .A(net3099),
    .Y(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[323] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2478),
    .C1(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2472),
    .A1(net2795),
    .Y(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[323]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[323] ),
    .B(net2948));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[323]_sg13g2_nor3_1_A  (.A(net1311),
    .B(net2795),
    .C(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[323]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[324] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net641),
    .C1(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2402),
    .A1(net2795),
    .Y(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2476),
    .B(net2472),
    .X(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[324] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y ),
    .A2(net2842),
    .Y(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[325] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net600),
    .C1(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2401),
    .A1(net2408),
    .Y(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2474));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2794),
    .B(net2906),
    .X(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[325] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[326]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2403),
    .B2(net786),
    .A2(net2899),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3278),
    .D(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[326] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2473));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[326]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[326]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[326] ),
    .B(net2950));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net963),
    .A2(net2472),
    .A1(net2285));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[327] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2898));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[327] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2403),
    .B2(net664),
    .A2(net2644),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[328] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[328] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y ),
    .A2(net2846),
    .Y(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y ),
    .A2(net3133));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2402),
    .B2(net733),
    .A2(net2686),
    .A1(net2795));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[329] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2400));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[329] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y ),
    .A2(net2842),
    .Y(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[329]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[329] ),
    .B(net2949));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1  (.B2(net3103),
    .C1(net2823),
    .B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[32] ),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2826));
 sg13g2_or2_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A  (.X(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X ),
    .B(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1  (.A2(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X ),
    .X(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_A_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1  (.B2(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X ),
    .B1(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ));
 sg13g2_nand2b_2 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N ),
    .A_N(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nor2b_2 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A  (.A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y ),
    .B_N(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N ),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y  (.B2(net3072),
    .C1(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ),
    .B1(net95),
    .A1(net2719),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N ),
    .A2(\i_snitch.consec_pc[0] ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(net2949),
    .B(net40),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2360),
    .B2(net861),
    .A2(net2904),
    .A1(net2767));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3257),
    .D(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[32] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2363));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[32] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y ),
    .A2(net2998),
    .Y(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net3027));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[330]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2405),
    .B2(net997),
    .A2(net2473),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[330] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2798),
    .B(net2693));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[330]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[330]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[330] ),
    .B(net2950));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[331]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2404),
    .B2(net709),
    .A2(net2680),
    .A1(net2797));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[331] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[331] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y ),
    .A2(net2845),
    .Y(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2403),
    .B2(net949),
    .A2(net2691),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3308),
    .D(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[332] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[332] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[268]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2846));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[332]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[332] ),
    .B(net2952));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2405),
    .B2(net976),
    .A2(net2689),
    .A1(net2798));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[333] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2474));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[333] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y ),
    .A2(net2843),
    .Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[333]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[333] ),
    .B(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2405),
    .B2(net947),
    .A2(net2687),
    .A1(net2798));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[334] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2474));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[334] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[302]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2844));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(net2958),
    .B(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[334]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[334]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[334] ),
    .B(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2404),
    .B2(net656),
    .A2(net2677),
    .A1(net2797));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[335] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[335] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y ),
    .A2(net2846),
    .Y(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y ),
    .A2(net3135));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3286),
    .D(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[336] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2473),
    .B2(net2263),
    .A2(net2668),
    .A1(net2798));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[336] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[272]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2843));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net451),
    .B(net2405));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[336]_sg13g2_nand2_1_A_1  (.Y(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_nand2_1_A_1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[336] ),
    .B(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2404),
    .B2(net723),
    .A2(net2663),
    .A1(net2797));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[337] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[337] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y ),
    .A2(net2845),
    .Y(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[337]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[337] ),
    .B(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2405),
    .B2(net672),
    .A2(net2473),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[338] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2798),
    .B(net2676));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[338] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[274]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_nand2_1_A_1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2844));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y ),
    .A2(net3129));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[339]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net1070),
    .A2(net2472),
    .A1(net2271));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[339] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2674));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[339]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[339]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[339] ),
    .B(net2947));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[161] ),
    .C1(net3027),
    .B1(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a21oi_1_A1_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[33] ),
    .Y(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2831));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[33] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2455),
    .B2(net2514),
    .A2(net2902),
    .A1(net2766));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net514),
    .B(net2359));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[33]_sg13g2_nand2_1_A_1  (.Y(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_nand2_1_A_1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[33] ),
    .B(net2825));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2403),
    .B2(net864),
    .A2(net2672),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3315),
    .D(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[340] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[340] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[276]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2845));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(net2959),
    .B(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[340]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[340]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[340] ),
    .B(net2952));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net948),
    .A2(net2472),
    .A1(net2269));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3264),
    .D(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[341] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2670));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[341] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y ),
    .A2(net2841),
    .Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[341] ),
    .B(net2948));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[309]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[342]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2403),
    .B2(net743),
    .A2(net2652),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[342] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[342] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[310]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2847));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[343]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2403),
    .B2(net891),
    .A2(net2647),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3308),
    .D(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[343] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2399));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[343] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y ),
    .A2(net2846),
    .Y(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2404),
    .B2(net879),
    .A2(net2666),
    .A1(net2797));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3315),
    .D(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[344] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2400),
    .A2(net310));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[344] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[280]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2845));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y ),
    .A2(net3137));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net781),
    .A2(net2472),
    .A1(net2267));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[345] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2662));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[345] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[345]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[345] ),
    .B(net2948));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2401),
    .B2(net703),
    .A2(net2472),
    .A1(net2255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[346] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2660));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[346] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y ),
    .A2(net3116));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net894),
    .A2(net2472),
    .A1(net2253));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[347] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2658));
 sg13g2_nor2b_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_nor2b_1_B_N  (.A(net3115),
    .B_N(\i_snitch.i_snitch_regfile.mem[347] ),
    .Y(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[347]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[347] ),
    .A2(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[348]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2401),
    .B2(net909),
    .A2(net2473),
    .A1(net2246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[348] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2794),
    .B(net2655));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[348]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[348]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[348] ),
    .B(net2950));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2405),
    .B2(net1073),
    .A2(net2473),
    .A1(net2251));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[349] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2798),
    .B(net2653));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[349] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[317]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2843));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1  (.B2(net3099),
    .C1(net2821),
    .B1(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[34] ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2824));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_and2_1_A_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1 ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_and2_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A  (.B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_A ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B ),
    .B2(net93),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C ),
    .A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B ));
 sg13g2_and3_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B_sg13g2_and3_1_X  (.X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B ),
    .A(net3033),
    .B(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_B ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ),
    .C1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_C_sg13g2_nand2_1_Y_B ));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1_sg13g2_nor4_1_Y  (.A(net3079),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ),
    .C(net96),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_nand4_1_A_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(net3076),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1 ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_nor3_1_C  (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_A ),
    .B(net76),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ));
 sg13g2_or4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_A_Y ),
    .B(net2744),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X ),
    .D(net95),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B  (.A(net2515),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B_Y ),
    .A(net2515),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y  (.A(net2848),
    .B(net52),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nand3_1_Y  (.B(net2926),
    .C(net2925),
    .A(net2922),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y  (.A(net2928),
    .B(net51),
    .C(net2848),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C  (.A(net2848),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ));
 sg13g2_or2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_or2_1_X  (.X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ),
    .B(net3081),
    .A(net3083));
 sg13g2_or3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1 ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B ),
    .C(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_Y_sg13g2_nand3_1_A_Y),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B_sg13g2_o21ai_1_Y  (.B1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_C1_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_B ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_A ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y ),
    .B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ),
    .B2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X ),
    .A2(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .A1(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C  (.B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y ),
    .A(net44),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B_sg13g2_inv_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_B ),
    .A(net92));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y  (.B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2 ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_C ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y  (.A(net96),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and4_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ));
 sg13g2_nor4_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A ));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A_C ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_B_sg13g2_nand4_1_Y_C ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_and2_1_X  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ),
    .B(net2815),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B ));
 sg13g2_or2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B  (.X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_C_sg13g2_nor2_1_Y_A ));
 sg13g2_nand2b_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ),
    .A_N(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_C1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y  (.A(net96),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_C ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ),
    .B(net93));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_nor3_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor4_1_A_C ));
 sg13g2_or3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A_sg13g2_or3_1_A  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_Y_A ),
    .B(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_A ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_D_B ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B ),
    .X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .B2(net2815),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_C_sg13g2_and2_1_X_B ),
    .A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D ),
    .A2(net2744),
    .A1(net2928));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1_sg13g2_nor4_1_Y  (.A(net3077),
    .B(net83),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_D_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1 ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ));
 sg13g2_and3_2 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C  (.X(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_X ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A_sg13g2_nand2b_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A ),
    .B(net3093),
    .A_N(net40));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ),
    .B1(net95),
    .B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .A2(net2719),
    .A1(\i_req_arb.data_i[37] ));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C  (.B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ),
    .C(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_A ),
    .A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2974),
    .B2(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3006),
    .A1(\i_snitch.i_snitch_regfile.mem[34] ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3224),
    .D(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[34] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2485),
    .C1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_nor3_1_A_Y ),
    .B1(net2454),
    .A1(net2765),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2912));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[34]_sg13g2_nor3_1_A  (.A(net1326),
    .B(net2765),
    .C(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_nor3_1_A_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2405),
    .B2(net964),
    .A2(net2473),
    .A1(net2245));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[350] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2798),
    .B(net2650));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[350] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y ),
    .A2(net2843),
    .Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[350]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[350] ),
    .B(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[351]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2403),
    .B2(net813),
    .A2(net2645),
    .A1(net2796));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[351] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[351]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2400));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[352]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[352] ),
    .A2(net3124),
    .Y(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2941));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[352]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2398),
    .B2(net957),
    .A2(net2904),
    .A1(net2880));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3255),
    .D(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[352] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[352]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2393));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[353] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2470),
    .B2(net2513),
    .A2(net2901),
    .A1(net2881));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net457),
    .B(net2395));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[353] ),
    .A2(net2951));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[289]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[354] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2485),
    .C1(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2471),
    .A1(net2879),
    .Y(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2912));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[354]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[354] ),
    .B(net3117));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[354]_sg13g2_nor3_1_A  (.A(net1334),
    .B(net2879),
    .C(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[354]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[354]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[354] ),
    .A2(net2801));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[355]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[355] ),
    .A2(net3121),
    .Y(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[355] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2478),
    .C1(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2471),
    .A1(net2879),
    .Y(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[355]_sg13g2_nor3_1_A  (.A(net1206),
    .B(net2879),
    .C(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[355]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[356] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2476),
    .C1(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2469),
    .A1(net2879),
    .Y(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[356]_sg13g2_nor3_1_A  (.A(net1284),
    .B(net2879),
    .C(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[356]_sg13g2_o21ai_1_A1  (.B1(net2969),
    .Y(\i_snitch.i_snitch_regfile.mem[356]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[356] ),
    .A2(net2803));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3222),
    .D(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[357] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2408),
    .C1(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2471),
    .A1(net2878),
    .Y(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2906));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[357]_sg13g2_nor3_1_A  (.A(net1337),
    .B(net2878),
    .C(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[357]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[357]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[357] ),
    .A2(net2801));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[358]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[358] ),
    .A2(net124),
    .Y(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[358]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net1102),
    .A2(net2899),
    .A1(net2881));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[358] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[358]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2470));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[359]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net1031),
    .A2(net2469),
    .A1(net2285));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[359] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2878),
    .B(net2898));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[359]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[359]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[359] ),
    .A2(net2800));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[35] ),
    .A2(net3006),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2979));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_mux2_1_A0_X ),
    .B2(net3101),
    .A2(net2824),
    .A1(\i_snitch.i_snitch_regfile.mem[35] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2933),
    .C1(\i_snitch.i_snitch_regfile.mem[131]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y ),
    .A1(net3089),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A1(net2637),
    .B1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1 ),
    .X(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1 ),
    .A1(net2931),
    .A2(net70));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1_sg13g2_o21ai_1_Y_B1 ),
    .B1(net95),
    .B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .A2(net2719),
    .A1(\i_req_arb.data_i[38] ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A1(net2637));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[35] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_nor3_1_A_Y ),
    .B1(net2454),
    .A1(net2765),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[35]_sg13g2_nor3_1_A  (.A(net1279),
    .B(net2764),
    .C(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_nor3_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[360]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[360] ),
    .A2(net3133),
    .Y(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[360]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net737),
    .A2(net2644),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[360] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[360]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[360]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[360] ),
    .A2(net2808));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[361]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[361] ),
    .A2(net3123),
    .Y(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2946));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[361]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2398),
    .B2(net795),
    .A2(net2686),
    .A1(net2880));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[361] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2393));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[361]_sg13g2_o21ai_1_A1  (.B1(net2969),
    .Y(\i_snitch.i_snitch_regfile.mem[361]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[361] ),
    .A2(net2802));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[362]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[362] ),
    .A2(net3132),
    .Y(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[362]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net930),
    .A2(net2470),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3270),
    .D(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[362] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[362]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2881),
    .B(net2693));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[363]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net848),
    .A2(net2680),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[363] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[363]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[363]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[363] ),
    .A2(net2807));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[364]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[364] ),
    .A2(net3134),
    .Y(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[364]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net839),
    .A2(net2691),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[364] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[364]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[364]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[364] ),
    .A2(net2808));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[365] ),
    .A2(net3130),
    .Y(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net1014),
    .A2(net2689),
    .A1(net2881));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3286),
    .D(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[365] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2470));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[365]_sg13g2_o21ai_1_A1  (.B1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[365]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[365] ),
    .A2(net2804));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[366] ),
    .A2(net3130),
    .Y(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2943));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net1194),
    .A2(net2687),
    .A1(net2881));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[366] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2471));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[366]_sg13g2_o21ai_1_A1  (.B1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[366]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[366] ),
    .A2(net2805));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[367]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[367] ),
    .A2(net3135),
    .Y(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[367]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net895),
    .A2(net2677),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3293),
    .D(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[367] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[367]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[367]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[367] ),
    .A2(net2808));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[368] ),
    .A2(net3129),
    .Y(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2943));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net1094),
    .A2(net2470),
    .A1(net2263));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3286),
    .D(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[368] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2881),
    .B(net2668));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[368]_sg13g2_o21ai_1_A1  (.B1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[368]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[368] ),
    .A2(net2805));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[369]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[369] ),
    .A2(net3135),
    .Y(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[369]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net888),
    .A2(net2663),
    .A1(net2883));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[369] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[369]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[369]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[369] ),
    .A2(net2807));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[36] ),
    .A2(net3008),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2980));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[100]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_mux2_1_A0_X ),
    .B2(net3103),
    .A2(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[36] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2933),
    .A2(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3224),
    .D(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[36] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2476),
    .C1(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_nor3_1_A_Y ),
    .B1(net2454),
    .A1(net2767),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[36]_sg13g2_nor3_1_A  (.A(net1379),
    .B(net2767),
    .C(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_nor3_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[370] ),
    .A2(net3129),
    .Y(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2943));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net986),
    .A2(net2470),
    .A1(net2272));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[370] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2881),
    .B(net2676));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[370]_sg13g2_o21ai_1_A1  (.B1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[370]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[370] ),
    .A2(net2805));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[371]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[371] ),
    .A2(net3116),
    .Y(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[371]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net988),
    .A2(net2469),
    .A1(net2271));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[371] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[371]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2878),
    .B(net2674));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[372]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[372] ),
    .A2(net3137),
    .Y(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[372]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net985),
    .A2(net2672),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3316),
    .D(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[372] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[372]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[372]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[372] ),
    .A2(net2806));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[373] ),
    .A2(net3119),
    .Y(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net1141),
    .A2(net2469),
    .A1(net2269));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[373] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2878),
    .B(net2670));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[373]_sg13g2_o21ai_1_A1  (.B1(net2969),
    .Y(\i_snitch.i_snitch_regfile.mem[373]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[373] ),
    .A2(net2802));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[374]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net753),
    .A2(net2652),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3314),
    .D(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[374] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[374]_sg13g2_o21ai_1_A1  (.B1(net2971),
    .Y(\i_snitch.i_snitch_regfile.mem[374]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[374] ),
    .A2(net2808));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[375]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2396),
    .B2(net904),
    .A2(net2647),
    .A1(net2882));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3310),
    .D(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[375] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2392));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[375]_sg13g2_o21ai_1_A1  (.B1(net2972),
    .Y(\i_snitch.i_snitch_regfile.mem[375]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[375] ),
    .A2(net2808));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[376]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[376] ),
    .A2(net3137),
    .Y(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[376]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2397),
    .B2(net1191),
    .A2(net2666),
    .A1(net2882));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[376] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2393),
    .A2(net310));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[376]_sg13g2_o21ai_1_A1  (.B1(net2972),
    .Y(\i_snitch.i_snitch_regfile.mem[376]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[376] ),
    .A2(net2806));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[377] ),
    .A2(net3119),
    .Y(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2941));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[377] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2469),
    .B2(net2267),
    .A2(net2662),
    .A1(net2878));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net467),
    .B(net2394));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[377]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[377]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[377] ),
    .A2(net2800));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[378] ),
    .A2(net3116),
    .Y(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net1021),
    .A2(net2469),
    .A1(net2255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3213),
    .D(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[378] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2878),
    .B(net2660));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[378]_sg13g2_o21ai_1_A1  (.B1(net2968),
    .Y(\i_snitch.i_snitch_regfile.mem[378]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[378] ),
    .A2(net2800));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[379] ),
    .A2(net3116),
    .Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net1000),
    .A2(net2469),
    .A1(net2253));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[379] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2878),
    .B(net2658));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[379] ),
    .B(net2800),
    .Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[347]_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[37] ),
    .A2(net2824),
    .Y(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2821));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_1  (.A1(\i_snitch.i_snitch_regfile.mem[37] ),
    .A2(net3001),
    .Y(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_a21oi_1_A1_1_Y ),
    .B1(net2974));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[37]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[37] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[37]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2408),
    .C1(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_nor3_1_A_Y ),
    .B1(net2455),
    .A1(net2765),
    .Y(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2906));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[37]_sg13g2_nor3_1_A  (.A(net1340),
    .B(net2765),
    .C(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[37]_sg13g2_nor3_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[380]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[380] ),
    .A2(net3126),
    .Y(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[380]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2394),
    .B2(net1173),
    .A2(net2469),
    .A1(net2246));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[380] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[380]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2884),
    .B(net2656));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[381]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2395),
    .B2(net1022),
    .A2(net2470),
    .A1(net2250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[381] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2881),
    .B(net2654));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[381]_sg13g2_o21ai_1_A1  (.B1(net2970),
    .Y(\i_snitch.i_snitch_regfile.mem[381]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[381] ),
    .A2(net2804));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[382] ),
    .A2(net3127),
    .Y(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2943));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2397),
    .B2(net1125),
    .A2(net2470),
    .A1(net2245));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[382] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2883),
    .B(net2650));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[382]_sg13g2_o21ai_1_A1  (.B1(net2972),
    .Y(\i_snitch.i_snitch_regfile.mem[382]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[382] ),
    .A2(net2804));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[383]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2394),
    .B2(net802),
    .A2(net2645),
    .A1(net2880));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3307),
    .D(\i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[383] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[383]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2393));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2388),
    .B2(net1077),
    .A2(net2903),
    .A1(net3039));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[384] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2386));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[384] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_inv_1_A_Y ),
    .A2(net3010));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0  (.S0(net3122),
    .A0(\i_snitch.i_snitch_regfile.mem[384] ),
    .A1(\i_snitch.i_snitch_regfile.mem[416] ),
    .A2(\i_snitch.i_snitch_regfile.mem[448] ),
    .A3(\i_snitch.i_snitch_regfile.mem[480] ),
    .S1(net3104),
    .X(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X_sg13g2_nand2_1_B_Y ),
    .A(net3093),
    .B(\i_snitch.i_snitch_regfile.mem[384]_sg13g2_mux4_1_A0_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3274),
    .D(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[385] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2514),
    .A2(net2902),
    .A1(net3040));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[385]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[385]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net495),
    .B(net2389));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[386] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2468),
    .A1(net3039),
    .Y(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0  (.S0(net3001),
    .A0(\i_snitch.i_snitch_regfile.mem[386] ),
    .A1(\i_snitch.i_snitch_regfile.mem[418] ),
    .A2(\i_snitch.i_snitch_regfile.mem[450] ),
    .A3(\i_snitch.i_snitch_regfile.mem[482] ),
    .S1(net2974),
    .X(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1  (.S0(net3117),
    .A0(\i_snitch.i_snitch_regfile.mem[386] ),
    .A1(\i_snitch.i_snitch_regfile.mem[418] ),
    .A2(\i_snitch.i_snitch_regfile.mem[450] ),
    .A3(\i_snitch.i_snitch_regfile.mem[482] ),
    .S1(net3102),
    .X(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1  (.B2(net3091),
    .C1(net2929),
    .B1(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_nand2_1_A_Y_sg13g2_nand3_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[386]_sg13g2_nor3_1_A  (.A(net1341),
    .B(net3039),
    .C(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[386]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[387] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net694),
    .C1(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2387),
    .A1(net3038),
    .Y(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2477),
    .B(net2466),
    .X(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[387] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y ),
    .A2(net3006));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0  (.S0(net3121),
    .A0(\i_snitch.i_snitch_regfile.mem[387] ),
    .A1(\i_snitch.i_snitch_regfile.mem[419] ),
    .A2(\i_snitch.i_snitch_regfile.mem[451] ),
    .A3(\i_snitch.i_snitch_regfile.mem[483] ),
    .S1(net3101),
    .X(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3092),
    .A2(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3219),
    .D(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[388] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net780),
    .C1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2388),
    .A1(net3039),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2475),
    .B(net2466),
    .X(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[388] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2919));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1  (.A1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_nand2b_2 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .A_N(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2b_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A  (.A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y ),
    .B_N(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .C1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ),
    .B1(net95),
    .A1(\i_req_arb.data_i[39] ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .A2(net2719));
 sg13g2_nor2b_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2b_1_Y  (.A(net40),
    .B_N(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2511),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0  (.S0(net3007),
    .A0(\i_snitch.i_snitch_regfile.mem[388] ),
    .A1(\i_snitch.i_snitch_regfile.mem[420] ),
    .A2(\i_snitch.i_snitch_regfile.mem[452] ),
    .A3(\i_snitch.i_snitch_regfile.mem[484] ),
    .S1(net2980),
    .X(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2957),
    .B1(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2962),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2640),
    .B(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[132]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1  (.A2(net2751),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .B1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[389] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2468),
    .A1(net674),
    .Y(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2387));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net3038),
    .B(net2905),
    .X(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[389] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2918));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0  (.S0(net3001),
    .A0(\i_snitch.i_snitch_regfile.mem[389] ),
    .A1(\i_snitch.i_snitch_regfile.mem[421] ),
    .A2(\i_snitch.i_snitch_regfile.mem[453] ),
    .A3(\i_snitch.i_snitch_regfile.mem[485] ),
    .S1(net2974),
    .X(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2640),
    .B(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[133]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1  (.A2(net2751),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ),
    .B1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[38] ),
    .A2(net2829),
    .Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2822));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[134]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[102]_sg13g2_o21ai_1_A1_Y ),
    .A1(net3088),
    .Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(net2637),
    .B2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net2719),
    .A1(\i_req_arb.data_i[41] ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A ),
    .A(net3086),
    .B(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_A ),
    .B(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1013),
    .A2(net2900),
    .A1(net2768));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3280),
    .D(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[38] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2456));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[38]_sg13g2_o21ai_1_A1  (.B1(net3013),
    .Y(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[38] ),
    .A2(net2990));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2389),
    .B2(net1145),
    .A2(net2899),
    .A1(net3040));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[390] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2467));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[390] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_inv_1_A_Y ),
    .A2(net3014));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0  (.S0(net124),
    .A0(\i_snitch.i_snitch_regfile.mem[390] ),
    .A1(\i_snitch.i_snitch_regfile.mem[422] ),
    .A2(\i_snitch.i_snitch_regfile.mem[454] ),
    .A3(\i_snitch.i_snitch_regfile.mem[486] ),
    .S1(net3107),
    .X(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3094),
    .A2(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[390]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2285),
    .A2(net2387),
    .A1(net1317));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3211),
    .D(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[391] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2897));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[391] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2918));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0  (.S0(net3001),
    .A0(\i_snitch.i_snitch_regfile.mem[391] ),
    .A1(\i_snitch.i_snitch_regfile.mem[423] ),
    .A2(\i_snitch.i_snitch_regfile.mem[455] ),
    .A3(\i_snitch.i_snitch_regfile.mem[487] ),
    .S1(net2974),
    .X(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[327]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[263]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2638),
    .B(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[135]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1  (.A2(net2751),
    .A1(net3084),
    .B1(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net760),
    .A2(net2644),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[392] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0  (.S0(net3133),
    .A0(\i_snitch.i_snitch_regfile.mem[392] ),
    .A1(\i_snitch.i_snitch_regfile.mem[424] ),
    .A2(\i_snitch.i_snitch_regfile.mem[456] ),
    .A3(\i_snitch.i_snitch_regfile.mem[488] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1  (.S0(net3019),
    .A0(\i_snitch.i_snitch_regfile.mem[392] ),
    .A1(\i_snitch.i_snitch_regfile.mem[424] ),
    .A2(\i_snitch.i_snitch_regfile.mem[456] ),
    .A3(\i_snitch.i_snitch_regfile.mem[488] ),
    .S1(net2990),
    .X(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2959),
    .B1(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2965),
    .Y(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1  (.Y(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X ),
    .B2(net3096),
    .A2(\i_snitch.i_snitch_regfile.mem[264]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[328]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2388),
    .B2(net800),
    .A2(net2685),
    .A1(net3039));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[393] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2386));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0  (.S0(net3123),
    .A0(\i_snitch.i_snitch_regfile.mem[393] ),
    .A1(\i_snitch.i_snitch_regfile.mem[425] ),
    .A2(\i_snitch.i_snitch_regfile.mem[457] ),
    .A3(\i_snitch.i_snitch_regfile.mem[489] ),
    .S1(net3103),
    .X(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1  (.S0(net3009),
    .A0(\i_snitch.i_snitch_regfile.mem[393] ),
    .A1(\i_snitch.i_snitch_regfile.mem[425] ),
    .A2(\i_snitch.i_snitch_regfile.mem[457] ),
    .A3(\i_snitch.i_snitch_regfile.mem[489] ),
    .S1(net2982),
    .X(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2  (.Y(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[329]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X ),
    .A1(net2967));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X ),
    .A1(net3093),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[394] ),
    .A2(net3027),
    .Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_a21o_1_A1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2468),
    .B2(net2283),
    .A2(net2389),
    .A1(net1251));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3274),
    .D(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[394] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3040),
    .B(net2694));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0  (.S0(net3121),
    .A0(\i_snitch.i_snitch_regfile.mem[394] ),
    .A1(\i_snitch.i_snitch_regfile.mem[426] ),
    .A2(\i_snitch.i_snitch_regfile.mem[458] ),
    .A3(\i_snitch.i_snitch_regfile.mem[490] ),
    .S1(net3110),
    .X(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3094),
    .A2(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[266]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A1(net3088),
    .B1(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ),
    .B(net2509),
    .Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .A(net3078),
    .B(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1  (.A2(net2722),
    .A1(\i_snitch.inst_addr_o[10] ),
    .B1(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2722),
    .A1(\i_snitch.inst_addr_o[10] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net883),
    .A2(net2680),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3316),
    .D(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[395] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0  (.S0(net3021),
    .A0(\i_snitch.i_snitch_regfile.mem[395] ),
    .A1(\i_snitch.i_snitch_regfile.mem[427] ),
    .A2(\i_snitch.i_snitch_regfile.mem[459] ),
    .A3(\i_snitch.i_snitch_regfile.mem[491] ),
    .S1(net2992),
    .X(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[331]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2958),
    .B1(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2965),
    .Y(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1  (.A2(net2753),
    .A1(net3133),
    .B1(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[395]_sg13g2_o21ai_1_A1  (.B1(net3097),
    .Y(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[395] ),
    .A2(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net1121),
    .A2(net2691),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[396] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0  (.S0(net3134),
    .A0(\i_snitch.i_snitch_regfile.mem[396] ),
    .A1(\i_snitch.i_snitch_regfile.mem[428] ),
    .A2(\i_snitch.i_snitch_regfile.mem[460] ),
    .A3(\i_snitch.i_snitch_regfile.mem[492] ),
    .S1(net3113),
    .X(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1  (.S0(net3024),
    .A0(\i_snitch.i_snitch_regfile.mem[396] ),
    .A1(\i_snitch.i_snitch_regfile.mem[428] ),
    .A2(\i_snitch.i_snitch_regfile.mem[460] ),
    .A3(\i_snitch.i_snitch_regfile.mem[492] ),
    .S1(net2991),
    .X(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2  (.A1(net2965),
    .A2(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[332]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X ),
    .A1(net3096),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[396]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2389),
    .B2(net850),
    .A2(net2689),
    .A1(net3040));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[397] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2467));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0  (.S0(net3130),
    .A0(\i_snitch.i_snitch_regfile.mem[397] ),
    .A1(\i_snitch.i_snitch_regfile.mem[429] ),
    .A2(\i_snitch.i_snitch_regfile.mem[461] ),
    .A3(\i_snitch.i_snitch_regfile.mem[493] ),
    .S1(net3109),
    .X(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1  (.S0(net3017),
    .A0(\i_snitch.i_snitch_regfile.mem[397] ),
    .A1(\i_snitch.i_snitch_regfile.mem[429] ),
    .A2(\i_snitch.i_snitch_regfile.mem[461] ),
    .A3(\i_snitch.i_snitch_regfile.mem[493] ),
    .S1(net2988),
    .X(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2  (.Y(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[333]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_1_X ),
    .A1(net2963));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X ),
    .A1(net3094),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[397]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2390),
    .B2(net1130),
    .A2(net2687),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3292),
    .D(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[398] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2468));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0  (.S0(net3130),
    .A0(\i_snitch.i_snitch_regfile.mem[398] ),
    .A1(\i_snitch.i_snitch_regfile.mem[430] ),
    .A2(\i_snitch.i_snitch_regfile.mem[462] ),
    .A3(\i_snitch.i_snitch_regfile.mem[494] ),
    .S1(net3109),
    .X(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X ),
    .A1(net3095),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[398]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[398] ),
    .B(net3028));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net793),
    .A2(net2677),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[399] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0  (.S0(net3135),
    .A0(\i_snitch.i_snitch_regfile.mem[399] ),
    .A1(\i_snitch.i_snitch_regfile.mem[431] ),
    .A2(\i_snitch.i_snitch_regfile.mem[463] ),
    .A3(\i_snitch.i_snitch_regfile.mem[495] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1  (.S0(net3020),
    .A0(\i_snitch.i_snitch_regfile.mem[399] ),
    .A1(\i_snitch.i_snitch_regfile.mem[431] ),
    .A2(\i_snitch.i_snitch_regfile.mem[463] ),
    .A3(\i_snitch.i_snitch_regfile.mem[495] ),
    .S1(net2992),
    .X(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2959),
    .B1(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2966),
    .Y(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1  (.Y(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X ),
    .B2(net3097),
    .A2(\i_snitch.i_snitch_regfile.mem[303]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[335]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[39] ),
    .A2(net2824),
    .Y(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2821));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net1053),
    .A2(net2454),
    .A1(net2285));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3215),
    .D(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[39] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2898));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[39]_sg13g2_o21ai_1_A1  (.B1(net3011),
    .Y(\i_snitch.i_snitch_regfile.mem[39]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[39] ),
    .A2(net2975));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2262),
    .A2(net2389),
    .A1(net1225));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[400] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3040),
    .B(net2667));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0  (.S0(net3129),
    .A0(\i_snitch.i_snitch_regfile.mem[400] ),
    .A1(\i_snitch.i_snitch_regfile.mem[432] ),
    .A2(\i_snitch.i_snitch_regfile.mem[464] ),
    .A3(\i_snitch.i_snitch_regfile.mem[496] ),
    .S1(net3108),
    .X(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1  (.S0(net3016),
    .A0(\i_snitch.i_snitch_regfile.mem[400] ),
    .A1(\i_snitch.i_snitch_regfile.mem[432] ),
    .A2(\i_snitch.i_snitch_regfile.mem[464] ),
    .A3(\i_snitch.i_snitch_regfile.mem[496] ),
    .S1(net2987),
    .X(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2  (.A1(net2963),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[336]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ),
    .A1(net2954),
    .B1(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2641),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_B1 ),
    .A(net2993),
    .B(net2725));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X ),
    .A1(net3095),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2391),
    .B2(net975),
    .A2(net2663),
    .A1(net3042));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[401] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0  (.S0(net3135),
    .A0(\i_snitch.i_snitch_regfile.mem[401] ),
    .A1(\i_snitch.i_snitch_regfile.mem[433] ),
    .A2(\i_snitch.i_snitch_regfile.mem[465] ),
    .A3(\i_snitch.i_snitch_regfile.mem[497] ),
    .S1(net3112),
    .X(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1  (.S0(net3020),
    .A0(\i_snitch.i_snitch_regfile.mem[401] ),
    .A1(\i_snitch.i_snitch_regfile.mem[433] ),
    .A2(\i_snitch.i_snitch_regfile.mem[465] ),
    .A3(\i_snitch.i_snitch_regfile.mem[497] ),
    .S1(net2992),
    .X(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[337]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2958),
    .B1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2963),
    .Y(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X ),
    .A1(net3094),
    .B1(net2930),
    .X(\i_snitch.i_snitch_regfile.mem[401]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2272),
    .A2(net2389),
    .A1(net1164));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3283),
    .D(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[402] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3040),
    .B(net2675));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0  (.S0(net3129),
    .A0(\i_snitch.i_snitch_regfile.mem[402] ),
    .A1(\i_snitch.i_snitch_regfile.mem[434] ),
    .A2(\i_snitch.i_snitch_regfile.mem[466] ),
    .A3(\i_snitch.i_snitch_regfile.mem[498] ),
    .S1(net3108),
    .X(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1  (.S0(net3016),
    .A0(\i_snitch.i_snitch_regfile.mem[402] ),
    .A1(\i_snitch.i_snitch_regfile.mem[434] ),
    .A2(\i_snitch.i_snitch_regfile.mem[466] ),
    .A3(\i_snitch.i_snitch_regfile.mem[498] ),
    .S1(net2987),
    .X(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2  (.A1(net2964),
    .A2(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1  (.Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[402]_sg13g2_mux4_1_A0_X ),
    .B2(net3095),
    .A2(\i_snitch.i_snitch_regfile.mem[306]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[338]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2270),
    .A2(net2387),
    .A1(net1371));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3208),
    .D(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[403] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2673));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[403] ),
    .A1(\i_snitch.i_snitch_regfile.mem[435] ),
    .A2(\i_snitch.i_snitch_regfile.mem[467] ),
    .A3(\i_snitch.i_snitch_regfile.mem[499] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3091),
    .A2(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[275]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[403]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[403] ),
    .B(net3026));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net1111),
    .A2(net2672),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[404] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0  (.S0(net3137),
    .A0(\i_snitch.i_snitch_regfile.mem[404] ),
    .A1(\i_snitch.i_snitch_regfile.mem[436] ),
    .A2(\i_snitch.i_snitch_regfile.mem[468] ),
    .A3(\i_snitch.i_snitch_regfile.mem[500] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X ),
    .A1(net3096),
    .B1(net2931),
    .X(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[404]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[404] ),
    .B(net3029));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2268),
    .A2(net2387),
    .A1(net1220));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[405] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2669));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0  (.S0(net3120),
    .A0(\i_snitch.i_snitch_regfile.mem[405] ),
    .A1(\i_snitch.i_snitch_regfile.mem[437] ),
    .A2(\i_snitch.i_snitch_regfile.mem[469] ),
    .A3(\i_snitch.i_snitch_regfile.mem[501] ),
    .S1(net3101),
    .X(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1  (.S0(net3005),
    .A0(\i_snitch.i_snitch_regfile.mem[405] ),
    .A1(\i_snitch.i_snitch_regfile.mem[437] ),
    .A2(\i_snitch.i_snitch_regfile.mem[469] ),
    .A3(\i_snitch.i_snitch_regfile.mem[501] ),
    .S1(net2978),
    .X(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[277]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2962),
    .Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3092),
    .A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[341]_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A1(net3089),
    .B1(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(net2631),
    .Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2723),
    .A1(\i_snitch.inst_addr_o[21] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[406]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[406] ),
    .A2(net3030),
    .Y(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2992));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[406]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2391),
    .B2(net1100),
    .A2(net2652),
    .A1(net3042));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3316),
    .D(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[406] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2386));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[406]_sg13g2_o21ai_1_A1  (.B1(net3097),
    .Y(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[406] ),
    .A2(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net898),
    .A2(net2647),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[407] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2385));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[407] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net110));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B  (.A(net2636),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1  (.A1(\i_snitch.inst_addr_o[23] ),
    .A2(net2722),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1  (.B2(net2631),
    .C1(net2565),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .A2(net2548));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B  (.A(net2631),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0  (.S0(net3024),
    .A0(\i_snitch.i_snitch_regfile.mem[407] ),
    .A1(\i_snitch.i_snitch_regfile.mem[439] ),
    .A2(\i_snitch.i_snitch_regfile.mem[471] ),
    .A3(\i_snitch.i_snitch_regfile.mem[503] ),
    .S1(net2991),
    .X(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[343]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2959),
    .B1(\i_snitch.i_snitch_regfile.mem[279]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2965),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B  (.A(net2641),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1  (.B2(net3088),
    .C1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y ),
    .B1(net2849),
    .A1(net3074),
    .Y(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(net2753));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[408] ),
    .A2(net3030),
    .Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2993));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2390),
    .B2(net827),
    .A2(net2665),
    .A1(net3041));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[408] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2385));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0  (.S0(net3137),
    .A0(\i_snitch.i_snitch_regfile.mem[408] ),
    .A1(\i_snitch.i_snitch_regfile.mem[440] ),
    .A2(\i_snitch.i_snitch_regfile.mem[472] ),
    .A3(\i_snitch.i_snitch_regfile.mem[504] ),
    .S1(net3111),
    .X(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1  (.Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X ),
    .B2(net3096),
    .A2(\i_snitch.i_snitch_regfile.mem[312]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ),
    .A1(net3088),
    .B1(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1  (.A2(net2722),
    .A1(\i_snitch.inst_addr_o[24] ),
    .B1(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2266),
    .A2(net2387),
    .A1(net1179));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[409] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2661));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0  (.S0(net3119),
    .A0(\i_snitch.i_snitch_regfile.mem[409] ),
    .A1(\i_snitch.i_snitch_regfile.mem[441] ),
    .A2(\i_snitch.i_snitch_regfile.mem[473] ),
    .A3(\i_snitch.i_snitch_regfile.mem[505] ),
    .S1(net3100),
    .X(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1  (.S0(net3004),
    .A0(\i_snitch.i_snitch_regfile.mem[409] ),
    .A1(\i_snitch.i_snitch_regfile.mem[441] ),
    .A2(\i_snitch.i_snitch_regfile.mem[473] ),
    .A3(\i_snitch.i_snitch_regfile.mem[505] ),
    .S1(net2977),
    .X(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[345]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X ),
    .A1(net3092),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[409]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[40] ),
    .A2(net2826),
    .Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2821));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[104]_sg13g2_o21ai_1_A1_Y ),
    .A1(net3090),
    .Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[392]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1 ),
    .B1(net2637),
    .A1(\i_req_arb.data_i[43] ),
    .Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net2722));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X  (.A(net3082),
    .B(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1 ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ),
    .B(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2360),
    .B2(net821),
    .A2(net2643),
    .A1(net2770));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[40] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2363));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[40]_sg13g2_o21ai_1_A1  (.B1(net3019),
    .Y(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[40] ),
    .A2(net2982));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2254),
    .A2(net2387),
    .A1(net1262));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[410] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2659));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[410] ),
    .A1(\i_snitch.i_snitch_regfile.mem[442] ),
    .A2(\i_snitch.i_snitch_regfile.mem[474] ),
    .A3(\i_snitch.i_snitch_regfile.mem[506] ),
    .S1(net3099),
    .X(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1  (.S0(net3000),
    .A0(\i_snitch.i_snitch_regfile.mem[410] ),
    .A1(\i_snitch.i_snitch_regfile.mem[442] ),
    .A2(\i_snitch.i_snitch_regfile.mem[474] ),
    .A3(\i_snitch.i_snitch_regfile.mem[506] ),
    .S1(net2976),
    .X(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1  (.B2(net3091),
    .C1(net2929),
    .B1(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[346]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[282]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2466),
    .B2(net2252),
    .A2(net2387),
    .A1(net1176));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[411] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3038),
    .B(net2657));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0  (.S0(net3115),
    .A0(\i_snitch.i_snitch_regfile.mem[411] ),
    .A1(\i_snitch.i_snitch_regfile.mem[443] ),
    .A2(\i_snitch.i_snitch_regfile.mem[475] ),
    .A3(\i_snitch.i_snitch_regfile.mem[507] ),
    .S1(net3098),
    .X(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1  (.S0(net2999),
    .A0(\i_snitch.i_snitch_regfile.mem[411] ),
    .A1(\i_snitch.i_snitch_regfile.mem[443] ),
    .A2(\i_snitch.i_snitch_regfile.mem[475] ),
    .A3(\i_snitch.i_snitch_regfile.mem[507] ),
    .S1(net2973),
    .X(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.i_snitch_regfile.mem[379]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ),
    .C1(net2956),
    .B1(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X ),
    .A1(net3091),
    .B1(net2929),
    .X(\i_snitch.i_snitch_regfile.mem[411]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2246),
    .A2(net2389),
    .A1(net1129));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[412] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3040),
    .B(net2655));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[412] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_inv_1_A_Y ),
    .A2(net3012));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0  (.S0(net3126),
    .A0(\i_snitch.i_snitch_regfile.mem[412] ),
    .A1(\i_snitch.i_snitch_regfile.mem[444] ),
    .A2(\i_snitch.i_snitch_regfile.mem[476] ),
    .A3(\i_snitch.i_snitch_regfile.mem[508] ),
    .S1(net3106),
    .X(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2  (.A1(net3094),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[316]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .A1(net3088),
    .B1(\i_snitch.i_snitch_regfile.mem[156]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ),
    .B(net2511),
    .Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2720),
    .A1(\i_snitch.inst_addr_o[28] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[413] ),
    .A2(net3028),
    .Y(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2985));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2251),
    .A2(net2389),
    .A1(net1308));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3270),
    .D(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[413] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3040),
    .B(net2654));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[413]_sg13g2_o21ai_1_A1  (.B1(net3094),
    .Y(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[413] ),
    .A2(net2814));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2467),
    .B2(net2244),
    .A2(net2391),
    .A1(net1155));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[414] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net3042),
    .B(net2649));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0  (.S0(net3126),
    .A0(\i_snitch.i_snitch_regfile.mem[414] ),
    .A1(\i_snitch.i_snitch_regfile.mem[446] ),
    .A2(\i_snitch.i_snitch_regfile.mem[478] ),
    .A3(\i_snitch.i_snitch_regfile.mem[510] ),
    .S1(net3106),
    .X(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X ));
 sg13g2_mux4_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1  (.S0(net3015),
    .A0(\i_snitch.i_snitch_regfile.mem[414] ),
    .A1(\i_snitch.i_snitch_regfile.mem[446] ),
    .A2(\i_snitch.i_snitch_regfile.mem[478] ),
    .A3(\i_snitch.i_snitch_regfile.mem[510] ),
    .S1(net2985),
    .X(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2  (.Y(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[350]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X ),
    .A1(net2964));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2  (.A2(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X ),
    .A1(net3095),
    .B1(net2930),
    .X(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_a22oi_1_B2_Y ),
    .B1(net2388),
    .B2(net597),
    .A2(net2646),
    .A1(net3039));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[415] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2386));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[415] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y ),
    .A2(net110),
    .Y(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net2937));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y ),
    .A2(net3009));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[416]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[416] ),
    .A2(net3010),
    .Y(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2981));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[416]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2384),
    .B2(net886),
    .A2(net2903),
    .A1(net2861));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[416] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[416]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2380));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[417]_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[385] ),
    .C1(net2936),
    .B1(net2920),
    .A1(\i_snitch.i_snitch_regfile.mem[417] ),
    .Y(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2825));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[417] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2513),
    .A2(net2901),
    .A1(net2862));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[417]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[417]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net524),
    .B(net2381));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3217),
    .D(\i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[418] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2465),
    .A1(net2865),
    .Y(\i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[418]_sg13g2_nor3_1_A  (.A(net1339),
    .B(net2865),
    .C(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[418]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[419]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[419] ),
    .A2(net3006),
    .Y(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2979));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[419] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2463),
    .A1(net2860),
    .Y(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[419]_sg13g2_nor3_1_A  (.A(net1301),
    .B(net2860),
    .C(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[419]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1  (.B2(net3103),
    .C1(net2823),
    .B1(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[41] ),
    .Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2826));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2360),
    .B2(net841),
    .A2(net2685),
    .A1(net2767));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[41] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2363));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[105]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[41] ),
    .A2(net2982));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_a21oi_1_A1_Y ),
    .C1(net2642),
    .B1(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y ),
    .A1(net2955),
    .Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[393]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[137]_sg13g2_mux4_1_A0_1_X_sg13g2_nand2b_1_A_N_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(net2753),
    .A1(net3080));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[420] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2463),
    .A1(net2865),
    .Y(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[420]_sg13g2_nor3_1_A  (.A(net1315),
    .B(net2861),
    .C(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1  (.B1(net3091),
    .Y(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[420] ),
    .A2(net2811));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_A2 ),
    .A(net2940),
    .B(net3120));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[421] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2465),
    .A1(net2860),
    .Y(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[421]_sg13g2_nor3_1_A  (.A(net1328),
    .B(net2860),
    .C(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[421]_sg13g2_o21ai_1_A1  (.B1(net3091),
    .Y(\i_snitch.i_snitch_regfile.mem[421]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[421] ),
    .A2(net2810));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[422]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[422] ),
    .A2(net3014),
    .Y(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2986));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[422]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2381),
    .B2(net1101),
    .A2(net2899),
    .A1(net2862));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[422] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[422]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2464));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[423]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2284),
    .A2(net2384),
    .A1(net1356));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[423] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2860),
    .B(net2897));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[423]_sg13g2_o21ai_1_A1  (.B1(net3091),
    .Y(\i_snitch.i_snitch_regfile.mem[423]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[423] ),
    .A2(net2810));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[424]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net816),
    .A2(net2644),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[424] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[424]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2379));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[425]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2384),
    .B2(net779),
    .A2(net2685),
    .A1(net2861));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[425] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[425]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2380));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[426]_sg13g2_a21o_1_A1  (.A2(net3013),
    .A1(\i_snitch.i_snitch_regfile.mem[426] ),
    .B1(net2979),
    .X(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_a21o_1_A1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[426]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2465),
    .B2(net2283),
    .A2(net2381),
    .A1(net1185));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[426] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[426]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2862),
    .B(net2694));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net1068),
    .A2(net2679),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[427] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2379));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[427] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2828));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[267]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2631),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2636),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1  (.A2(net2722),
    .A1(\i_snitch.inst_addr_o[11] ),
    .B1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2722),
    .A1(\i_snitch.inst_addr_o[11] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1  (.A1(net2569),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(net90));
 sg13g2_nand3_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2_sg13g2_nand3_1_C  (.B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .C(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_A2 ),
    .A(net2569),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C  (.A(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B ),
    .C(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B ),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A  (.B(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1  (.B1(net90),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net2567),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor3_1_C  (.A(net2567),
    .B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .C(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor3_1_C_B ));
 sg13g2_and3_1 \i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C  (.X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_B ),
    .C(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[428]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net936),
    .A2(net2692),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[428] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[428]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2379));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[429]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2381),
    .B2(net805),
    .A2(net2689),
    .A1(net2862));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[429] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[429]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2464));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[42] ),
    .A2(net2827),
    .Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2822));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1168),
    .A2(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y ),
    .A1(net2282));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[42] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2768),
    .B(net2693));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[42] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_nand2_1_A_Y ),
    .B2(net3028),
    .A2(net2997),
    .A1(\i_snitch.i_snitch_regfile.mem[42]_sg13g2_inv_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[430]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[430] ),
    .A2(net3018),
    .Y(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2988));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[430] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2465),
    .B2(net2274),
    .A2(net2687),
    .A1(net2862));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[430]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net455),
    .B(net2381));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[431]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net829),
    .A2(net2677),
    .A1(net2864));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[431] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[431]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2379));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[432] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2262),
    .A2(net2667),
    .A1(net2862));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[432]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[432]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net438),
    .B(net2381));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[433]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net792),
    .A2(net2663),
    .A1(net2864));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[433] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[433]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2379));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[434]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2273),
    .A2(net2383),
    .A1(net1146));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[434] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[434]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2864),
    .B(net2675));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[435]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[435] ),
    .A2(net2999),
    .Y(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2973));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[435]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2270),
    .A2(net2384),
    .A1(net1255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[435] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2860),
    .B(net2673));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[436]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[436] ),
    .A2(net3023),
    .Y(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2993));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[436]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net1034),
    .A2(net2671),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[436] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2379));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[437]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2268),
    .A2(net2384),
    .A1(net1296));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[437] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[437]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2861),
    .B(net2669));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net801),
    .A2(net2651),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[438] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2379));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[438] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2829));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[278]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2510),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2632),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2635),
    .A2(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.A1(\i_snitch.inst_addr_o[22] ),
    .A2(net2723),
    .Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[438]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[438] ),
    .B(net3020));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[439]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2383),
    .B2(net757),
    .A2(net2647),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[439] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2379));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[439]_sg13g2_o21ai_1_A1  (.B1(net3096),
    .Y(\i_snitch.i_snitch_regfile.mem[439]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[439] ),
    .A2(net2812));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1  (.B2(net3112),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[43] ),
    .Y(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2828));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[139]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2361),
    .B2(net1079),
    .A2(net2680),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[43] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2281),
    .A2(net2363));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[43]_sg13g2_o21ai_1_A1  (.B1(net3021),
    .Y(\i_snitch.i_snitch_regfile.mem[43]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[43] ),
    .A2(net2994));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[440]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2383),
    .B2(net796),
    .A2(net2665),
    .A1(net2863));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[440] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2380));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[440]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[440] ),
    .B(net3022));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[441]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2266),
    .A2(net2384),
    .A1(net1186));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[441] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[441]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2861),
    .B(net2661));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[442] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2254),
    .A2(net2659),
    .A1(net2860));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[442]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[442]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net510),
    .B(net2384));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[443]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2463),
    .B2(net2252),
    .A2(net2384),
    .A1(net1285));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3210),
    .D(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[443] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[443]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2860),
    .B(net2657));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[444]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[444] ),
    .A2(net3012),
    .Y(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2985));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[444]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2246),
    .A2(net2381),
    .A1(net1202));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[444] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[444]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2862),
    .B(net2655));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2250),
    .A2(net2381),
    .A1(net1214));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[445] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2862),
    .B(net2653));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[445] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2827));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[285]_sg13g2_mux4_1_A0_X_sg13g2_a21o_1_A2_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .B(net2508),
    .Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(net2636),
    .A2(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2720),
    .A1(\i_snitch.inst_addr_o[29] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_A2  (.A1(net2695),
    .A2(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2540));
 sg13g2_inv_2 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[445]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[445] ),
    .B(net3015));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[446] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2464),
    .B2(net2244),
    .A2(net2649),
    .A1(net2864));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[446]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[446]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net454),
    .B(net2383));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[447]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[447] ),
    .A2(net3009),
    .Y(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2983));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[447]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2382),
    .B2(net933),
    .A2(net2646),
    .A1(net2863));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3305),
    .D(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[447] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2380));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[447]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[415]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[447] ),
    .A2(net2812));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[448]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2372),
    .B2(net742),
    .A2(net2903),
    .A1(net2739));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[448] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2378));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[448]_sg13g2_o21ai_1_A1  (.B1(net2962),
    .Y(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[448] ),
    .A2(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3279),
    .D(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[449] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2461),
    .B2(net2513),
    .A2(net2901),
    .A1(net2741));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net485),
    .B(net2373));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_o21ai_1_A1  (.B1(net3107),
    .Y(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[449] ),
    .A2(net3128));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[449]_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_B1 ),
    .A(\i_snitch.i_snitch_regfile.mem[449]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_mux2_1_A0_X ),
    .B2(net3113),
    .A2(net2829),
    .A1(\i_snitch.i_snitch_regfile.mem[44] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2934),
    .A2(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[140]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net1082),
    .A2(net2692),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3310),
    .D(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[44] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2277),
    .A2(net2363));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[44] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_nand2_1_A_Y ),
    .B2(net3029),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[44]_sg13g2_inv_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[450] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2462),
    .A1(net2739),
    .Y(\i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[450]_sg13g2_nor3_1_A  (.A(net1270),
    .B(net2739),
    .C(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[450]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3274),
    .D(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[451] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net675),
    .C1(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2372),
    .A1(net2738),
    .Y(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1_sg13g2_and2_1_X  (.A(net2478),
    .B(net2460),
    .X(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[451] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y ),
    .A2(net2841),
    .Y(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[452] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2460),
    .A1(net2739),
    .Y(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[452]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[452] ),
    .B(net2947));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[452]_sg13g2_nor3_1_A  (.A(net1281),
    .B(net2739),
    .C(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[452]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[453] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2462),
    .A1(net2738),
    .Y(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[453]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[453] ),
    .B(net2947));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[453]_sg13g2_nor3_1_A  (.A(net1321),
    .B(net2738),
    .C(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[453]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net856),
    .A2(net2899),
    .A1(net2742));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[454] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2461));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[454] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y ),
    .A2(net2843),
    .Y(\i_snitch.i_snitch_regfile.mem[454]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[455]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net1008),
    .A2(net2460),
    .A1(net2284));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[455] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2738),
    .B(net2897));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[455]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[455]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[455] ),
    .B(net2947));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[456]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net815),
    .A2(net2644),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3280),
    .D(\i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[456] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[456]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2377));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[457]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2376),
    .B2(net788),
    .A2(net2685),
    .A1(net2740));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[457] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[457]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2378));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3274),
    .D(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[458] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2462),
    .B2(net2283),
    .A2(net2694),
    .A1(net2742));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[458]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net513),
    .B(net2374));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[458]_sg13g2_o21ai_1_A1  (.B1(net2962),
    .Y(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[458] ),
    .A2(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[459]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net892),
    .A2(net2679),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[459] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2377));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[459]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[459]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[459] ),
    .B(net2953));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_mux2_1_A0_X ),
    .B2(net3108),
    .A2(net2830),
    .A1(\i_snitch.i_snitch_regfile.mem[45] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2934),
    .A2(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1046),
    .A2(net2690),
    .A1(net2768));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[45] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2456));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[45] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[45]_sg13g2_inv_1_A_Y ),
    .A2(net3031));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[460]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net762),
    .A2(net2691),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[460] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[460]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2377));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[461]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net1044),
    .A2(net2689),
    .A1(net2742));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[461] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[461]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2461));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2373),
    .B2(net1096),
    .A2(net2687),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[462] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2462));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[462] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[430]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[398]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[462]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2844));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[463]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net744),
    .A2(net2677),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3294),
    .D(\i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[463] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[463]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2377));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[464]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net983),
    .A2(net2461),
    .A1(net2262));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[464] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[464]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2742),
    .B(net2667));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[465]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net774),
    .A2(net2663),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[465] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[465]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2288),
    .A2(net2377));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[466]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net1123),
    .A2(net2461),
    .A1(net2273));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[466] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[466]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2742),
    .B(net2675));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net1159),
    .A2(net2460),
    .A1(net2270));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[467] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2738),
    .B(net2673));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[467] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[435]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[467]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2840));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[468]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2373),
    .B2(net905),
    .A2(net2671),
    .A1(net2741));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[468] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2377));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[468] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[436]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[404]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[468]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2845));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[469]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net943),
    .A2(net2460),
    .A1(net2268));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3262),
    .D(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[469] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[469]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2740),
    .B(net2669));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1  (.B2(net3109),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[46] ),
    .Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2830));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1124),
    .A2(net2687),
    .A1(net2768));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[46] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2456));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[46]_sg13g2_o21ai_1_A1  (.B1(net3017),
    .Y(\i_snitch.i_snitch_regfile.mem[46]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[46] ),
    .A2(net2988));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2375),
    .B2(net881),
    .A2(net2651),
    .A1(net2743));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[470] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2377));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[470] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[406]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2846));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(net2959),
    .B(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[342]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[470]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[470]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[470] ),
    .B(net2952));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[471]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2375),
    .B2(net716),
    .A2(net2647),
    .A1(net2743));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[471] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2377));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[471]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[471]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[471] ),
    .B(net2952));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2375),
    .B2(net862),
    .A2(net2665),
    .A1(net2743));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[472] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2378));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[472] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[440]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2845));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(net2959),
    .B(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[344]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[472]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[473]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net838),
    .A2(net2460),
    .A1(net2266));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[473] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[473]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2738),
    .B(net2661));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[474]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net1099),
    .A2(net2460),
    .A1(net2255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[474] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[474]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2738),
    .B(net2659));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[475]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2372),
    .B2(net826),
    .A2(net2460),
    .A1(net2252));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[475] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[475]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2738),
    .B(net2657));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net1120),
    .A2(net2461),
    .A1(net2247));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3267),
    .D(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[476] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2742),
    .B(net2656));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[476] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y ),
    .A2(net2841),
    .Y(\i_snitch.i_snitch_regfile.mem[476]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net932),
    .A2(net2461),
    .A1(net2250));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[477] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2742),
    .B(net2653));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[477] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[413]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_o21ai_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .A2(net2843));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B  (.A(net2958),
    .B(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[349]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[477]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[477]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[477] ),
    .B(net2950));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[478]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2374),
    .B2(net935),
    .A2(net2461),
    .A1(net2244));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[478] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[478]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2742),
    .B(net2649));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[479] ),
    .A2(net2949),
    .Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_a21o_1_A1_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[287]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[447]_sg13g2_o21ai_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2376),
    .B2(net789),
    .A2(net2645),
    .A1(net2740));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[479] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2378));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1  (.B1(net2967),
    .Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[479] ),
    .A2(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_A2 ),
    .A(net3026),
    .B(net2974));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[47] ),
    .A2(net2828),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2823));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y ),
    .C1(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[111]_sg13g2_o21ai_1_A1_Y ),
    .A1(net3090),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[399]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(net2637),
    .B2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net2725),
    .A1(\i_snitch.inst_addr_o[15] ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B  (.A(net2631),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D  (.B(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y ),
    .A(net2569),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y ));
 sg13g2_nand4_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C  (.B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A ),
    .C(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D ));
 sg13g2_or2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A_sg13g2_or2_1_X  (.X(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_A ),
    .B(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A(net2566));
 sg13g2_or2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D_sg13g2_or2_1_X  (.X(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_D ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ),
    .A(net2566));
 sg13g2_nor3_2 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C  (.A(net34),
    .B(net48),
    .C(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_and4_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y_sg13g2_and4_1_C  (.A(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .D(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ));
 sg13g2_nor4_2 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C  (.A(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .B(net48),
    .C(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y ),
    .D(net34));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B  (.A(net2566),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B ),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y  (.B1(net2567),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_xnor2_1_A_B ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ),
    .A1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .A(net2631),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_A2  (.B1(net2542),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net845),
    .A2(net2678),
    .A1(net2769));
 sg13g2_dfrbpq_2 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3299),
    .D(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[47] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2363));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[47]_sg13g2_o21ai_1_A1  (.B1(net3023),
    .Y(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[47] ),
    .A2(net2994));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[480]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2367),
    .B2(net973),
    .A2(net2903),
    .A1(net2855));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[480] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2521),
    .A2(net2366));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[480] ),
    .B(net2802),
    .Y(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[448]_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[480]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[481] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2514),
    .A2(net2902),
    .A1(net2857));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[481]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net447),
    .B(net2368));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[481]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[481] ),
    .A2(net2950));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[482] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2484),
    .C1(\i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2459),
    .A1(net2855),
    .Y(\i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2911));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[482]_sg13g2_nor3_1_A  (.A(net1307),
    .B(net2855),
    .C(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[482]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[483] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2478),
    .C1(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2457),
    .A1(net2856),
    .Y(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2910));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[483]_sg13g2_nor3_1_A  (.A(net1277),
    .B(net2854),
    .C(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[483]_sg13g2_o21ai_1_A1  (.B1(net2962),
    .Y(\i_snitch.i_snitch_regfile.mem[483]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[483] ),
    .A2(net2801));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[484]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[484] ),
    .A2(net3122),
    .Y(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2946));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[484] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2475),
    .C1(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2457),
    .A1(net2855),
    .Y(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2907));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[484]_sg13g2_nor3_1_A  (.A(net1313),
    .B(net2855),
    .C(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[484]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[485]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[485] ),
    .A2(net3117),
    .Y(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3218),
    .D(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[485] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2407),
    .C1(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2459),
    .A1(net2854),
    .Y(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2905));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[485]_sg13g2_nor3_1_A  (.A(net1249),
    .B(net2854),
    .C(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[485]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[486]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2369),
    .B2(net878),
    .A2(net2900),
    .A1(net2858));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3291),
    .D(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[486] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2286),
    .B(net2458));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[486]_sg13g2_o21ai_1_A1  (.B1(net2964),
    .Y(\i_snitch.i_snitch_regfile.mem[486]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[486] ),
    .A2(net2804));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[487]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[487] ),
    .A2(net3117),
    .Y(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[487]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2284),
    .A2(net2367),
    .A1(net1314));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[487] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[487]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2854),
    .B(net2897));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[488]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net882),
    .A2(net2644),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3280),
    .D(\i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[488] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[488]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2279),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[489]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2367),
    .B2(net875),
    .A2(net2685),
    .A1(net2855));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3275),
    .D(\i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[489] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[489]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2299),
    .A2(net2366));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1  (.B2(net3108),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[48] ),
    .Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2827));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[144]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1198),
    .A2(net2456),
    .A1(net2262));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[48] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2768),
    .B(net2667));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[48]_sg13g2_o21ai_1_A1  (.B1(net3018),
    .Y(\i_snitch.i_snitch_regfile.mem[48]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[48] ),
    .A2(net2987));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2459),
    .B2(net2283),
    .A2(net2369),
    .A1(net1241));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3277),
    .D(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[490] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2858),
    .B(net2694));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[490] ),
    .B(net2801),
    .Y(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B  (.A(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_a21oi_1_A1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[458]_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[490]_sg13g2_nor2_1_A_Y_sg13g2_nor3_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[491]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[491] ),
    .A2(net3135),
    .Y(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2945));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[491]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net1025),
    .A2(net2679),
    .A1(net2859));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[491] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[491]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[492]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net1112),
    .A2(net2691),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[492] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[492]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[493]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2369),
    .B2(net1017),
    .A2(net2690),
    .A1(net2858));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[493] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[493]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2290),
    .B(net2458));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[494]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2368),
    .B2(net952),
    .A2(net2688),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[494] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2275),
    .B(net2459));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[494]_sg13g2_o21ai_1_A1  (.B1(net2964),
    .Y(\i_snitch.i_snitch_regfile.mem[494]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[494] ),
    .A2(net2804));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[495]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net1001),
    .A2(net2678),
    .A1(net2859));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[495] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[495]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2264),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[496]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2262),
    .A2(net2369),
    .A1(net1248));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[496] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[496]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2858),
    .B(net2667));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[497]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net956),
    .A2(net2664),
    .A1(net2859));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[497] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[497]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[498]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2273),
    .A2(net2369),
    .A1(net1261));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3290),
    .D(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[498] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[498]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2858),
    .B(net2675));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[499]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2271),
    .A2(net2367),
    .A1(net1325));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[499] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2854),
    .B(net2674));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[499]_sg13g2_o21ai_1_A1  (.B1(net2961),
    .Y(\i_snitch.i_snitch_regfile.mem[499]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[499] ),
    .A2(net2800));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1  (.B2(net3109),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[49] ),
    .Y(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2830));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net1057),
    .A2(net2664),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[49] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2363));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[49]_sg13g2_o21ai_1_A1  (.B1(net3017),
    .Y(\i_snitch.i_snitch_regfile.mem[49]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[49] ),
    .A2(net2988));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[500]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2370),
    .B2(net969),
    .A2(net2671),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[500] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2260),
    .A2(net2365));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[500]_sg13g2_o21ai_1_A1  (.B1(net2965),
    .Y(\i_snitch.i_snitch_regfile.mem[500]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[500] ),
    .A2(net2806));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[501]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2268),
    .A2(net2367),
    .A1(net1189));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3263),
    .D(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[501] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[501]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2856),
    .B(net2669));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[502]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[502] ),
    .A2(net3135),
    .Y(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[502]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2368),
    .B2(net1109),
    .A2(net2651),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3321),
    .D(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[502] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2258),
    .A2(net2365));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[502]_sg13g2_o21ai_1_A1  (.B1(net2965),
    .Y(\i_snitch.i_snitch_regfile.mem[502]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[502] ),
    .A2(net2806));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[503]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[503] ),
    .A2(net3137),
    .Y(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[503]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2370),
    .B2(net784),
    .A2(net2647),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3318),
    .D(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[503] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[503]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2248),
    .A2(net2365));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[504]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2370),
    .B2(net868),
    .A2(net2665),
    .A1(net2857));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[504] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2366));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[504]_sg13g2_o21ai_1_A1  (.B1(net2966),
    .Y(\i_snitch.i_snitch_regfile.mem[504]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[504] ),
    .A2(net2806));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[505]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2266),
    .A2(net2367),
    .A1(net1199));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3212),
    .D(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[505] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[505]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2854),
    .B(net2661));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[506]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2254),
    .A2(net2367),
    .A1(net1136));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3206),
    .D(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[506] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[506]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2854),
    .B(net2659));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[507]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2457),
    .B2(net2253),
    .A2(net2367),
    .A1(net1222));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3209),
    .D(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[507] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[507]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2854),
    .B(net2658));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[508]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2247),
    .A2(net2369),
    .A1(net1324));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[508] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2858),
    .B(net2656));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[508]_sg13g2_o21ai_1_A1  (.B1(net2963),
    .Y(\i_snitch.i_snitch_regfile.mem[508]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[508] ),
    .A2(net2801));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[509] ),
    .A2(net3127),
    .Y(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2250),
    .A2(net2369),
    .A1(net1267));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3268),
    .D(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[509] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2858),
    .B(net2653));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[509]_sg13g2_o21ai_1_A1  (.B1(net2963),
    .Y(\i_snitch.i_snitch_regfile.mem[509]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[509] ),
    .A2(net2804));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_mux2_1_A0_X ),
    .B2(net3108),
    .A2(net2827),
    .A1(\i_snitch.i_snitch_regfile.mem[50] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1076),
    .A2(net2456),
    .A1(net2273));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3286),
    .D(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[50] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2768),
    .B(net2676));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[50] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_nand2_1_A_Y ),
    .B2(net3031),
    .A2(net2997),
    .A1(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_inv_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3284),
    .D(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[510] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2458),
    .B2(net2244),
    .A2(net2649),
    .A1(net2858));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[510]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[510]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net453),
    .B(net2369));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_a21o_1_A1  (.A2(net3123),
    .A1(\i_snitch.i_snitch_regfile.mem[511] ),
    .B1(net2941),
    .X(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_a21o_1_A1_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2371),
    .B2(net842),
    .A2(net2645),
    .A1(net2856));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[511] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2242),
    .A2(net2366));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[511] ),
    .B(net2802),
    .Y(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[479]_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[511]_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_mux2_1_A0_X ),
    .B2(net3100),
    .A2(net2824),
    .A1(\i_snitch.i_snitch_regfile.mem[51] ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2933),
    .C1(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y ),
    .A1(net3089),
    .Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[403]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(net2723),
    .A1(\i_snitch.inst_addr_o[19] ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .A(net2631),
    .B(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net978),
    .A2(net2454),
    .A1(net2271));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[51] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2674));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[51] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_nand2_1_A_Y ),
    .B2(net3026),
    .A2(net2998),
    .A1(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_inv_1_A_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_mux2_1_A0_X ),
    .B2(net3114),
    .A2(net2828),
    .A1(\i_snitch.i_snitch_regfile.mem[52] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_1  (.Y(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_1_Y ),
    .B1(net2994),
    .B2(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3022),
    .A1(\i_snitch.i_snitch_regfile.mem[52] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2934),
    .A2(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net880),
    .A2(net2672),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[52] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[52]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2364));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[53] ),
    .A2(net2825),
    .Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2821));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2978),
    .B2(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3004),
    .A1(\i_snitch.i_snitch_regfile.mem[53] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[117]_sg13g2_nor2_1_A_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net867),
    .A2(net2455),
    .A1(net2269));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[53] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2670));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_mux2_1_A0_X ),
    .B2(net3112),
    .A2(net2828),
    .A1(\i_snitch.i_snitch_regfile.mem[54] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_1  (.Y(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_1_Y ),
    .B1(net2992),
    .B2(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3021),
    .A1(\i_snitch.i_snitch_regfile.mem[54] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2934),
    .A2(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net1117),
    .A2(net2652),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3320),
    .D(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[54] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[54]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2364));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_mux2_1_A0_X ),
    .B2(net3111),
    .A2(net2829),
    .A1(\i_snitch.i_snitch_regfile.mem[55] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_1  (.Y(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_1_Y ),
    .B1(net2994),
    .B2(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3022),
    .A1(\i_snitch.i_snitch_regfile.mem[55] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2934),
    .A2(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[151]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net1352),
    .A2(net2648),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[55] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[55]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2364));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[56] ),
    .A2(net2828),
    .Y(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2823));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2993),
    .B2(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3023),
    .A1(\i_snitch.i_snitch_regfile.mem[56] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2833),
    .Y(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[120]_sg13g2_nor2_1_A_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2362),
    .B2(net920),
    .A2(net2665),
    .A1(net2769));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[56] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[56]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2256),
    .A2(net2364));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1  (.B2(net3100),
    .C1(net2821),
    .B1(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[57] ),
    .Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2824));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net830),
    .A2(net2454),
    .A1(net2267));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3215),
    .D(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[57] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2662));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[57]_sg13g2_o21ai_1_A1  (.B1(net3004),
    .Y(\i_snitch.i_snitch_regfile.mem[57]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[57] ),
    .A2(net2977));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1  (.B2(net3100),
    .C1(net2821),
    .B1(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[58] ),
    .Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2824));
 sg13g2_or3_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C  (.A(\i_snitch.i_snitch_regfile.mem[410]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_B1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X ),
    .B(net2509),
    .Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2  (.B1(net2633),
    .Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y ),
    .A1(net2634),
    .A2(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2720),
    .A1(\i_snitch.inst_addr_o[26] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net981),
    .A2(net2454),
    .A1(net2255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[58] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2660));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[58]_sg13g2_o21ai_1_A1  (.B1(net3004),
    .Y(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[58] ),
    .A2(net2977));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_mux2_1_A0_X ),
    .B2(net3100),
    .A2(net2824),
    .A1(\i_snitch.i_snitch_regfile.mem[59] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_1  (.Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_1_Y ),
    .B1(net2977),
    .B2(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3004),
    .A1(\i_snitch.i_snitch_regfile.mem[59] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.A1(net2933),
    .A2(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net1071),
    .A2(net2454),
    .A1(net2253));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[59] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[59]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2764),
    .B(net2658));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[60] ),
    .A2(net2826),
    .Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2821));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y ),
    .B1(net2977),
    .B2(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3012),
    .A1(\i_snitch.i_snitch_regfile.mem[60] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2  (.B1(net2832),
    .Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[124]_sg13g2_nor2_1_A_1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_A1_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2359),
    .B2(net1011),
    .A2(net2455),
    .A1(net2247));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3269),
    .D(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[60] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[60]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2766),
    .B(net2656));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1  (.B2(net3106),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[61] ),
    .Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2827));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2360),
    .B2(net923),
    .A2(net2456),
    .A1(net2251));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3270),
    .D(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[61] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2768),
    .B(net2654));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[61]_sg13g2_o21ai_1_A1  (.B1(net3012),
    .Y(\i_snitch.i_snitch_regfile.mem[61]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[61] ),
    .A2(net2985));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1  (.B2(net3106),
    .C1(net2822),
    .B1(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_mux2_1_A0_X ),
    .A1(\i_snitch.i_snitch_regfile.mem[62] ),
    .Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2827));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_X_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_a221oi_1_A1_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2361),
    .B2(net1040),
    .A2(net2456),
    .A1(net2245));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[62] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2768),
    .B(net2650));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[126]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[62] ),
    .A2(net2986));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1  (.Y(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[62]_sg13g2_o21ai_1_A1_Y ),
    .B2(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[414]_sg13g2_mux4_1_A0_1_X_sg13g2_a22oi_1_A2_Y ),
    .A1(net2954));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_mux2_1_A0_X ),
    .B2(net3103),
    .A2(net2826),
    .A1(\i_snitch.i_snitch_regfile.mem[63] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_1  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_1_Y ),
    .B1(net2983),
    .B2(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_nand2b_1_A_N_Y ),
    .A2(net3009),
    .A1(\i_snitch.i_snitch_regfile.mem[63] ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y ),
    .A1(net2933));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2  (.B2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .C1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ),
    .B1(net2637),
    .A1(\i_snitch.inst_addr_o[31] ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(net2720));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S  (.A0(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0 ),
    .A1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B ),
    .S(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X ));
 sg13g2_a21o_2 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1  (.A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0 ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1 ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ),
    .B(net2549),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X ));
 sg13g2_nand2_2 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ),
    .B(net2549));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1  (.A1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A2 ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0 ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0 ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N ),
    .A1(net3145),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B ));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y_sg13g2_nor4_1_D  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y_sg13g2_nand3_1_C_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B_X ),
    .D(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_B ));
 sg13g2_or3_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B_sg13g2_or3_1_X  (.A(net96),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_B ),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_A_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nand3_1_C_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B  (.B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_A ),
    .A(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_xnor2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xnor2_1_B  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X ));
 sg13g2_xor2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B  (.B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y ),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X ));
 sg13g2_a21o_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X_sg13g2_a21o_1_B1  (.A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_A2_1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_B ));
 sg13g2_xnor2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y  (.A1(net2570),
    .A2(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y ),
    .A_N(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2b_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A  (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y ),
    .B_N(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A_Y ));
 sg13g2_and2_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B(net2512),
    .X(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_and2_1_A_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2360),
    .B2(net812),
    .A2(net2646),
    .A1(net2767));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[63] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2363));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1  (.B2(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .C1(net2834),
    .B1(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_nand2b_1_A_N_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[64] ),
    .Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2842));
 sg13g2_nor4_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C  (.A(net2642),
    .B(\i_snitch.i_snitch_regfile.mem[256]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y ),
    .D(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y ));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_A2 ),
    .A1(net3009));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .A2(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A1(net2700));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .B(net2602),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2354),
    .B2(net765),
    .A2(net2904),
    .A1(net2785));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3257),
    .D(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[64] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[64]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[64] ),
    .A1(\i_snitch.i_snitch_regfile.mem[96] ),
    .S(net3124),
    .X(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_mux2_1_A0_X ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[65] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2452),
    .B2(net2514),
    .A2(net2902),
    .A1(net2784));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[65] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_Y ),
    .B2(net2979),
    .A2(net2842),
    .A1(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_inv_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net458),
    .B(net2353));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[65] ),
    .B(net3120),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[33]_sg13g2_nand2_1_A_1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_1_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1  (.B2(net2933),
    .C1(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[353]_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_A1_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .A2(net3088));
 sg13g2_a21oi_2 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1  (.B1(net35),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net112),
    .A1(net113));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .A_N(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2b_2 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A  (.A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .B_N(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y  (.B2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ),
    .C1(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ),
    .B1(net95),
    .A1(\i_snitch.inst_addr_o[1] ),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N ),
    .A2(net2719));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(net2941),
    .B(net40),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_B_N_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A  (.A(net36),
    .B(net2509),
    .Y(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[66]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[66] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[66]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2485),
    .C1(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_nor3_1_A_Y ),
    .B1(net2451),
    .A1(net2783),
    .Y(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2912));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[66]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[66] ),
    .A1(\i_snitch.i_snitch_regfile.mem[98] ),
    .S(net3117),
    .X(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[66]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3026),
    .A_N(\i_snitch.i_snitch_regfile.mem[66] ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[66]_sg13g2_nor3_1_A  (.A(net1333),
    .B(net2783),
    .C(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[66]_sg13g2_nor3_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[67]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[67] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[67]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_nor3_1_A_Y ),
    .B1(net2451),
    .A1(net2782),
    .Y(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[67]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[67] ),
    .A1(\i_snitch.i_snitch_regfile.mem[99] ),
    .S(net3120),
    .X(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[67]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3026),
    .A_N(\i_snitch.i_snitch_regfile.mem[67] ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[67]_sg13g2_nor3_1_A  (.A(net1219),
    .B(net2782),
    .C(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_nor3_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[68]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3224),
    .D(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[68] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[68]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2476),
    .C1(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_nor3_1_A_Y ),
    .B1(net2452),
    .A1(net2784),
    .Y(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2908));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[68]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[68] ),
    .A1(\i_snitch.i_snitch_regfile.mem[100] ),
    .S(net3123),
    .X(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[68]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3032),
    .A_N(\i_snitch.i_snitch_regfile.mem[68] ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[68]_sg13g2_nor3_1_A  (.A(net1237),
    .B(net2784),
    .C(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[68]_sg13g2_nor3_1_A_Y ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[69]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[69] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[69]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2408),
    .C1(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_nor3_1_A_Y ),
    .B1(net2451),
    .A1(net2782),
    .Y(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2906));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[69]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3026),
    .A_N(\i_snitch.i_snitch_regfile.mem[69] ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[69]_sg13g2_nor3_1_A  (.A(net1288),
    .B(net2782),
    .C(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_nor3_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[69]_sg13g2_o21ai_1_A1  (.B1(net3099),
    .Y(\i_snitch.i_snitch_regfile.mem[69]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[69] ),
    .A2(net3117));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[70] ),
    .A2(net2846),
    .Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net1103),
    .A2(net2900),
    .A1(net2786));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3280),
    .D(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[70] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2287),
    .B(net2453));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[70] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y ),
    .A2(net2950),
    .Y(\i_snitch.i_snitch_regfile.mem[70]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net2942));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[71] ),
    .A2(net2841),
    .Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net987),
    .A2(net2451),
    .A1(net2285));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[71] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2782),
    .B(net2898));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[71] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y ),
    .A2(net2947),
    .Y(\i_snitch.i_snitch_regfile.mem[71]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net2940));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[72] ),
    .A2(net2842),
    .Y(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2354),
    .B2(net900),
    .A2(net2643),
    .A1(net2785));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3303),
    .D(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[72] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2278),
    .A2(net2357));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[72] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y ),
    .A2(net2952),
    .Y(\i_snitch.i_snitch_regfile.mem[72]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net2944));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[73]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[73] ),
    .A2(net2842),
    .Y(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[73]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2354),
    .B2(net794),
    .A2(net2686),
    .A1(net2785));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3302),
    .D(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[73] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2300),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[73]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[73] ),
    .A1(\i_snitch.i_snitch_regfile.mem[105] ),
    .S(net3123),
    .X(\i_snitch.i_snitch_regfile.mem[73]_sg13g2_mux2_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net919),
    .A2(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .A1(net2283));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3270),
    .D(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[74] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2786),
    .B(net2694));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[74] ),
    .B(net2995));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[74]_sg13g2_o21ai_1_A1  (.B1(net3110),
    .Y(\i_snitch.i_snitch_regfile.mem[74]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[74] ),
    .A2(net3132));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[75]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[75] ),
    .A2(net2846),
    .Y(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[75]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net934),
    .A2(net2679),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3319),
    .D(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[75] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2280),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[75]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[75] ),
    .A1(\i_snitch.i_snitch_regfile.mem[107] ),
    .S(net3136),
    .X(\i_snitch.i_snitch_regfile.mem[75]_sg13g2_mux2_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[76]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2354),
    .B2(net814),
    .A2(net2691),
    .A1(net2785));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3310),
    .D(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[76] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2276),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[76]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[76] ),
    .A1(\i_snitch.i_snitch_regfile.mem[108] ),
    .S(net3133),
    .X(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[76]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[76]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[76] ),
    .B(net2991));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net1115),
    .A2(net2690),
    .A1(net2786));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3295),
    .D(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[77] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2291),
    .B(net2453));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[77] ),
    .A1(\i_snitch.i_snitch_regfile.mem[109] ),
    .S(net3131),
    .X(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_mux2_1_A0_X ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[77]_sg13g2_o21ai_1_A1  (.B1(net2988),
    .Y(\i_snitch.i_snitch_regfile.mem[77]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[77] ),
    .A2(net3017));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[78] ),
    .A2(net2844),
    .Y(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net1091),
    .A2(net2688),
    .A1(net2786));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3296),
    .D(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[78] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2274),
    .B(net2453));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[78]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[78] ),
    .A1(\i_snitch.i_snitch_regfile.mem[110] ),
    .S(net3130),
    .X(\i_snitch.i_snitch_regfile.mem[78]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[79] ),
    .A2(net2845),
    .Y(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net977),
    .A2(net2678),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3297),
    .D(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[79] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2265),
    .A2(net2357));
 sg13g2_inv_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[79] ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y ),
    .A2(net2953),
    .Y(\i_snitch.i_snitch_regfile.mem[79]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(net2945));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[80] ),
    .A2(net2844),
    .Y(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3288),
    .D(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[80] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2453),
    .B2(net2262),
    .A2(net2667),
    .A1(net2786));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[80] ),
    .A1(\i_snitch.i_snitch_regfile.mem[112] ),
    .S(net3131),
    .X(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[80]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[80]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net523),
    .B(net2355));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[81]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[81] ),
    .A2(net2845),
    .Y(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[81]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2355),
    .B2(net1203),
    .A2(net2664),
    .A1(net2786));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3298),
    .D(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[81] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2289),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[81]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[81] ),
    .A1(\i_snitch.i_snitch_regfile.mem[113] ),
    .S(net3130),
    .X(\i_snitch.i_snitch_regfile.mem[81]_sg13g2_mux2_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net1010),
    .A2(net2453),
    .A1(net2273));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[82] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2786),
    .B(net2676));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[82] ),
    .A1(\i_snitch.i_snitch_regfile.mem[114] ),
    .S(net3129),
    .X(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[82]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[82]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[82] ),
    .B(net2987));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net929),
    .A2(net2451),
    .A1(net2271));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[83] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2783),
    .B(net2674));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[83] ),
    .A1(\i_snitch.i_snitch_regfile.mem[115] ),
    .S(net3120),
    .X(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[83]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[83]_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[83] ),
    .B(net2977));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[84]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net994),
    .A2(net2672),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3322),
    .D(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[84] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2261),
    .A2(net2358));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[84]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[84] ),
    .A1(\i_snitch.i_snitch_regfile.mem[116] ),
    .S(net3138),
    .X(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[84]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[84]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3030),
    .A_N(\i_snitch.i_snitch_regfile.mem[84] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net877),
    .A2(net2452),
    .A1(net2269));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[85] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2783),
    .B(net2670));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3027),
    .A_N(\i_snitch.i_snitch_regfile.mem[85] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[85]_sg13g2_o21ai_1_A1  (.B1(net3100),
    .Y(\i_snitch.i_snitch_regfile.mem[85]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[85] ),
    .A2(net3120));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[86]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net769),
    .A2(net2652),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3320),
    .D(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[86] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2259),
    .A2(net2358));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[86]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[86] ),
    .A1(\i_snitch.i_snitch_regfile.mem[118] ),
    .S(net3136),
    .X(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[86]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[86]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3029),
    .A_N(\i_snitch.i_snitch_regfile.mem[86] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[87]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net939),
    .A2(net2648),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3323),
    .D(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[87] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2249),
    .A2(net2358));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[87]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[87] ),
    .A1(\i_snitch.i_snitch_regfile.mem[119] ),
    .S(net3138),
    .X(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[87]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[87]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3030),
    .A_N(\i_snitch.i_snitch_regfile.mem[87] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[88]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2356),
    .B2(net766),
    .A2(net2666),
    .A1(net2787));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3324),
    .D(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[88] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2358),
    .A2(net2257));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[88]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3030),
    .A_N(\i_snitch.i_snitch_regfile.mem[88] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[88]_sg13g2_o21ai_1_A1  (.B1(net3111),
    .Y(\i_snitch.i_snitch_regfile.mem[88]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[88] ),
    .A2(net3138));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[89] ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net962),
    .A2(net2451),
    .A1(net2267));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3215),
    .D(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[89] ),
    .CLK(clknet_leaf_113_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2782),
    .B(net2662));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[89]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[89] ),
    .A1(\i_snitch.i_snitch_regfile.mem[121] ),
    .S(net3119),
    .X(\i_snitch.i_snitch_regfile.mem[89]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[90] ),
    .A2(net2840),
    .Y(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2834));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net1110),
    .A2(net2451),
    .A1(net2255));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3214),
    .D(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[90] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2782),
    .B(net2660));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[90]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[90] ),
    .A1(\i_snitch.i_snitch_regfile.mem[122] ),
    .S(net3119),
    .X(\i_snitch.i_snitch_regfile.mem[90]_sg13g2_mux2_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net1038),
    .A2(net2451),
    .A1(net2253));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3265),
    .D(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[91] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2783),
    .B(net2658));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[91] ),
    .A1(\i_snitch.i_snitch_regfile.mem[123] ),
    .S(net3119),
    .X(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[91]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[91]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3027),
    .A_N(\i_snitch.i_snitch_regfile.mem[91] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2353),
    .B2(net1037),
    .A2(net2452),
    .A1(net2247));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3266),
    .D(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[92] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2784),
    .B(net2656));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3026),
    .A_N(\i_snitch.i_snitch_regfile.mem[92] ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[92]_sg13g2_o21ai_1_A1  (.B1(net3100),
    .Y(\i_snitch.i_snitch_regfile.mem[92]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[92] ),
    .A2(net3126));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[93] ),
    .A2(net2843),
    .Y(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2354),
    .B2(net1131),
    .A2(net2453),
    .A1(net2251));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3270),
    .D(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[93] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2784),
    .B(net2654));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[93]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[93] ),
    .A1(\i_snitch.i_snitch_regfile.mem[125] ),
    .S(net3126),
    .X(\i_snitch.i_snitch_regfile.mem[93]_sg13g2_mux2_1_A0_X ));
 sg13g2_a21oi_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1  (.A1(\i_snitch.i_snitch_regfile.mem[94] ),
    .A2(net2843),
    .Y(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_Y ),
    .B1(net2835));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2355),
    .B2(net876),
    .A2(net2453),
    .A1(net2245));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3285),
    .D(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[94] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net2786),
    .B(net2650));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[94]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[94] ),
    .A1(\i_snitch.i_snitch_regfile.mem[126] ),
    .S(net3127),
    .X(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_mux2_1_A0_X ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[95]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2354),
    .B2(net731),
    .A2(net2646),
    .A1(net2785));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3304),
    .D(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[95] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2243),
    .A2(net2357));
 sg13g2_mux2_1 \i_snitch.i_snitch_regfile.mem[95]_sg13g2_mux2_1_A0  (.A0(\i_snitch.i_snitch_regfile.mem[95] ),
    .A1(\i_snitch.i_snitch_regfile.mem[127] ),
    .S(net3124),
    .X(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_mux2_1_A0_X ));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[95]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[95]_sg13g2_nand2b_1_A_N_Y ),
    .B(net3027),
    .A_N(\i_snitch.i_snitch_regfile.mem[95] ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[96]_sg13g2_a22oi_1_B2  (.Y(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2410),
    .B2(net872),
    .A2(net2904),
    .A1(net2869));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3257),
    .D(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[96] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D ),
    .A1(net2522),
    .A2(net2413));
 sg13g2_nand2b_1 \i_snitch.i_snitch_regfile.mem[96]_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_nand2b_1_A_N_Y ),
    .B(net2983),
    .A_N(\i_snitch.i_snitch_regfile.mem[96] ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3276),
    .D(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[97] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .B1(net2449),
    .B2(net2514),
    .A2(net2902),
    .A1(net2868));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_nand2_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_A ),
    .A(net494),
    .B(net2409));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1  (.B1(net2832),
    .Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[97] ),
    .A2(net3026));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_1  (.B1(net3101),
    .Y(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[97] ),
    .A2(net2951));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3221),
    .D(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[98] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2485),
    .C1(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_Y ),
    .B1(net2449),
    .A1(net2867),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2912));
 sg13g2_nor2_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A  (.A(\i_snitch.i_snitch_regfile.mem[98] ),
    .B(net2800),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_B ),
    .A(net3016),
    .B(net2989));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1  (.B1(net2831),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a22oi_1_A1_Y ));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A  (.A(net1358),
    .B(net2868),
    .C(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_Y ));
 sg13g2_nand2b_2 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nand2b_1_B  (.Y(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .B(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .A_N(net2867));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B  (.A(net2867),
    .B(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_2 \i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_Y  (.A(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ),
    .B(net2506),
    .Y(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ));
 sg13g2_dfrbpq_1 \i_snitch.i_snitch_regfile.mem[99]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3273),
    .D(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.i_snitch_regfile.mem[99] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_a221oi_1 \i_snitch.i_snitch_regfile.mem[99]_sg13g2_dfrbpq_1_Q_D_sg13g2_a221oi_1_Y  (.B2(net2477),
    .C1(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_nor3_1_A_Y ),
    .B1(net2448),
    .A1(net2866),
    .Y(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_dfrbpq_1_Q_D ),
    .A2(net2909));
 sg13g2_nor3_1 \i_snitch.i_snitch_regfile.mem[99]_sg13g2_nor3_1_A  (.A(net1364),
    .B(net2866),
    .C(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_nor3_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.i_snitch_regfile.mem[99]_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[67]_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_snitch.i_snitch_regfile.mem[99]_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.i_snitch_regfile.mem[99] ),
    .A2(net2801));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[10] ),
    .Q(\i_snitch.inst_addr_o[10] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3313),
    .D(\i_snitch.pc_d[11] ),
    .Q(\i_snitch.inst_addr_o[11] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3328),
    .D(\i_snitch.pc_d[12] ),
    .Q(\i_snitch.inst_addr_o[12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.pc_d[13] ),
    .Q(\i_snitch.inst_addr_o[13] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_xnor2_1 \i_snitch.inst_addr_o[13]_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ),
    .A(\i_snitch.inst_addr_o[13] ),
    .B(net2528));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[14] ),
    .Q(\i_snitch.inst_addr_o[14] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[15] ),
    .Q(\i_snitch.inst_addr_o[15] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[16] ),
    .Q(\i_snitch.inst_addr_o[16] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3317),
    .D(\i_snitch.pc_d[17] ),
    .Q(\i_snitch.inst_addr_o[17] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_a21o_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1  (.A2(net2528),
    .A1(\i_snitch.inst_addr_o[18] ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1 ),
    .X(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X ));
 sg13g2_a21oi_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1  (.A1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1_A1 ),
    .A2(net41),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1 ));
 sg13g2_and2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1_sg13g2_and2_1_X  (.A(\i_snitch.inst_addr_o[17] ),
    .B(net2528),
    .X(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1 ));
 sg13g2_a21o_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1  (.A2(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2 ),
    .A1(net41),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X ),
    .X(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X_sg13g2_a21oi_1_A2  (.A1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A2(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A  (.Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B ));
 sg13g2_and2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_and2_1_B  (.A(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2 ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B ),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nor3_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y  (.A(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B ));
 sg13g2_nor2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.inst_addr_o[19] ),
    .B(net2525),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A ));
 sg13g2_and2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B_sg13g2_and2_1_X  (.A(\i_snitch.inst_addr_o[19] ),
    .B(net2525),
    .X(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1  (.A1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y ),
    .A2(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_nand2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_B1 ),
    .A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_nand2b_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1 ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N_B ),
    .A_N(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_nand2_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B ));
 sg13g2_o21ai_1 \i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B_sg13g2_o21ai_1_Y  (.B1(net2525),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_B ),
    .A1(\i_snitch.inst_addr_o[19] ),
    .A2(\i_snitch.inst_addr_o[20] ));
 sg13g2_a221oi_1 \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1  (.B2(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2 ),
    .C1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y ),
    .A1(\i_snitch.inst_addr_o[18] ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ),
    .A2(net2724));
 sg13g2_a221oi_1 \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y  (.B2(net2934),
    .C1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[50]_sg13g2_a22oi_1_A1_Y ),
    .A1(net3088),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2 ),
    .A2(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_and2_1 \i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A  (.A(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2 ),
    .B(net2512),
    .X(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_and2_1_A_X ));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[18] ),
    .Q(\i_snitch.inst_addr_o[18] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_inv_2 \i_snitch.inst_addr_o[18]_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1355));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.pc_d[19] ),
    .Q(\i_snitch.inst_addr_o[19] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3256),
    .D(\i_snitch.pc_d[1] ),
    .Q(\i_snitch.inst_addr_o[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3309),
    .D(\i_snitch.pc_d[20] ),
    .Q(\i_snitch.inst_addr_o[20] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[21] ),
    .Q(\i_snitch.inst_addr_o[21] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3327),
    .D(\i_snitch.pc_d[22] ),
    .Q(\i_snitch.inst_addr_o[22] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[23] ),
    .Q(\i_snitch.inst_addr_o[23] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3313),
    .D(\i_snitch.pc_d[24] ),
    .Q(\i_snitch.inst_addr_o[24] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[25] ),
    .Q(\i_snitch.inst_addr_o[25] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[26] ),
    .Q(\i_snitch.inst_addr_o[26] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[27] ),
    .Q(\i_snitch.inst_addr_o[27] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3305),
    .D(\i_snitch.pc_d[28] ),
    .Q(\i_snitch.inst_addr_o[28] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[29] ),
    .Q(\i_snitch.inst_addr_o[29] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[30] ),
    .Q(\i_snitch.inst_addr_o[30] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 \i_snitch.inst_addr_o[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3312),
    .D(\i_snitch.pc_d[31] ),
    .Q(\i_snitch.inst_addr_o[31] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_nand2_1 \i_snitch.pc_d[0]_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[0] ),
    .A(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A ),
    .C(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.consec_pc[0] ),
    .Y(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y ));
 sg13g2_nand4_1 \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nand4_1_A  (.B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ),
    .C(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_Y ),
    .A(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_nand3_1_B_Y ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_C ),
    .D(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y  (.B1(net1174),
    .Y(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_A ),
    .A1(net2302),
    .A2(net2518));
 sg13g2_nand3_1 \i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y  (.B(net49),
    .C(net2312),
    .A(net2751),
    .Y(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[10] ),
    .A1(net2305),
    .A2(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2520),
    .A2(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2760),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .A2(net2626));
 sg13g2_xnor2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2b_2 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ),
    .A_N(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B  (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .C(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_C ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2717),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y  (.A1(net2706),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A ),
    .B1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2610),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .C1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2547),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2543),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .A2(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor3_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B(net33),
    .C(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C ),
    .Y(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_A_C ),
    .A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2552),
    .A2(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[394]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(net2684),
    .A1(net2745),
    .S(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .X(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand3_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C  (.B(net2313),
    .C(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.inst_addr_o[10] ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[10] ),
    .B(net2306),
    .C(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_B1 ),
    .A(net990),
    .B(net2306));
 sg13g2_a21o_1 \i_snitch.pc_d[11]_sg13g2_a21o_1_A2  (.A2(\i_snitch.pc_d[11] ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1 ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_B1 ),
    .X(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X ));
 sg13g2_nor4_2 \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A  (.A(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_D ),
    .B(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C_Y ),
    .C(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_C ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y ),
    .D(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X ));
 sg13g2_nand4_1 \i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C  (.B(\i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1_Y ),
    .C(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C_Y ),
    .D(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B_X ));
 sg13g2_a22oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[11] ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2307),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_2 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1 ),
    .A(net1385));
 sg13g2_xnor2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1 ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B ));
 sg13g2_and2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B_sg13g2_and2_1_X  (.A(net3072),
    .B(net2536),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1 ),
    .C(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2 ),
    .A(\i_snitch.inst_addr_o[11] ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y  (.B(net414),
    .C(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .A(net2519),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C  (.B(net414),
    .C(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .A(net2762),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B  (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A_Y ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y ),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B_X ));
 sg13g2_or3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X  (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B ),
    .C(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C ),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C ));
 sg13g2_nor3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ),
    .C(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B ));
 sg13g2_a21oi_2 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2 ),
    .A1(net45));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B_Y ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y  (.B(net3078),
    .C(net2537),
    .A(\i_snitch.inst_addr_o[10] ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net3078),
    .A2(net2537),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.inst_addr_o[10] ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_A2_Y ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_C ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2759),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2307));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B(net2629));
 sg13g2_nand3_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A ),
    .A1(net2541),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_inv_2 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1 ),
    .A(net2696));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1 ),
    .A2(net2579));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_B1 ),
    .A(net2748),
    .B(net2579));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2749),
    .B(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2546));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2572),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2588),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A(net2586),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2581),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(net2577));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2596),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2558),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2558),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2596),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2552),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2715),
    .A2(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2706),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2572),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2538));
 sg13g2_o21ai_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2584),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2594),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net2557),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_or2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A(net2580));
 sg13g2_nor2_1 \i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2610),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[12] ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2308),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_2 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1 ),
    .A(net1400));
 sg13g2_xnor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1 ),
    .B(net2527));
 sg13g2_and2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1 ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2 ),
    .X(\i_snitch.pc_d[12]_sg13g2_mux2_1_A1_A0 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2519),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_or2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A  (.X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2  (.B2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ),
    .C1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A_Y ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1 ),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_Y ),
    .A2(net2759));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B  (.A(net2763),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B_Y ));
 sg13g2_or2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1 ),
    .A(net2759));
 sg13g2_or3_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X  (.A(net2853),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B_sg13g2_a221oi_1_C1  (.B2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ),
    .C1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_B ),
    .B1(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_B_sg13g2_nor3_1_B_Y ),
    .Y(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C ),
    .A2(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y  (.B1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_B2_sg13g2_or3_1_C_X ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C ),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1_sg13g2_and2_1_X  (.A(net3144),
    .B(net3142),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or3_1_X_C_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_nor2b_2 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2_sg13g2_nor2b_1_Y  (.A(net3073),
    .B_N(net3148),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B2 ));
 sg13g2_and3_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A ),
    .A(\i_snitch.inst_addr_o[11] ),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_B ));
 sg13g2_or2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A  (.X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B_sg13g2_nor2_1_Y  (.A(\i_snitch.inst_addr_o[12] ),
    .B(net2527),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_C ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_X_A_sg13g2_or2_1_A_X_sg13g2_nand3_1_B_A ),
    .A(\i_snitch.inst_addr_o[12] ),
    .B(net2527));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y  (.A(net2309),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2717),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2706),
    .C1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2614),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_xnor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .A(net101),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_and4_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D  (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .C(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C ),
    .D(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X ));
 sg13g2_inv_2 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A ));
 sg13g2_xor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A ));
 sg13g2_xor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X  (.B(net55),
    .A(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y ),
    .A2(net33));
 sg13g2_a21oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_Y ),
    .A1(net67),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2b_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2572),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .B1(net2538));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2580),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2599),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2561),
    .B(net123),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1_Y ),
    .A1(net2709),
    .A2(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2561),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2561),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2580),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2597),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .S(net88),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_and2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2592),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y ),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B ),
    .A1(net2745),
    .A2(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2696),
    .B(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A  (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B(net2626),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_A_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[12]_sg13g2_mux2_1_A1  (.A0(\i_snitch.pc_d[12]_sg13g2_mux2_1_A1_A0 ),
    .A1(\i_snitch.pc_d[12] ),
    .S(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_A1 ),
    .X(\i_snitch.pc_d[12]_sg13g2_mux2_1_A1_X ));
 sg13g2_a21o_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X  (.A2(net2305),
    .A1(net1375),
    .B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[13] ));
 sg13g2_a221oi_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1  (.B2(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2 ),
    .C1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C_Y ),
    .B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1 ),
    .A1(\i_req_arb.data_i[43] ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A_X ));
 sg13g2_inv_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2 ),
    .A(\i_snitch.inst_addr_o[13] ));
 sg13g2_and2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X  (.A(net2313),
    .B(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C  (.A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_a221oi_1_B1_B2 ),
    .B(net2305),
    .C(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .A1(net2718),
    .A2(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y  (.A1(net73),
    .A2(net2851),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B ));
 sg13g2_or2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .A(net2717));
 sg13g2_nor2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A  (.A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .B(net2626),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor2_1_A_Y ));
 sg13g2_nor4_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ),
    .C(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .D(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2551),
    .A2(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2749),
    .A2(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2684),
    .B(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ));
 sg13g2_a21oi_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2697),
    .A2(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_B ),
    .B1(net2541));
 sg13g2_o21ai_1 \i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D ),
    .A1(net2610),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2309),
    .Y(\i_snitch.pc_d[14] ),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1363));
 sg13g2_a221oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2761),
    .C1(net2308),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2519),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2762),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[14] ),
    .B(net2527));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.inst_addr_o[13] ),
    .B(net2528));
 sg13g2_a22oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2629),
    .A2(net2851),
    .A1(net74));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand4_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .C(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y ),
    .D(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A ),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X  (.B(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y  (.A(net2566),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_X_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B ));
 sg13g2_and2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A ),
    .A1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_inv_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y_A1 ),
    .A(net46));
 sg13g2_nand3b_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y  (.B(net46),
    .C(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B ),
    .A_N(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C ),
    .A(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B ));
 sg13g2_nor4_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B  (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y ),
    .C(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .D(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y ));
 sg13g2_nand3_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y_sg13g2_nand3_1_A  (.B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .C(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A_Y ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_Y_sg13g2_nor4_1_B_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_C ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A2  (.A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B_Y ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_C1 ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_or2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y  (.A(net2567),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ));
 sg13g2_nor3_2 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .B(net48),
    .C(net34),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .A(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xnor2_1_B  (.Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[269]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(net55),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A1(net2566),
    .A2(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y  (.A(net67),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1  (.B2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A_X ),
    .C1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_C1 ),
    .B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y ),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X ));
 sg13g2_and2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .A1(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y_A ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2706),
    .C1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2546),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2697),
    .A2(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_A2 ),
    .B1(net2541));
 sg13g2_a21o_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(net2551),
    .B1(\i_snitch.i_snitch_regfile.mem[270]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(net2749),
    .A2(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2684),
    .B(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_B1 ),
    .B(\i_snitch.inst_addr_o[14] ),
    .A_N(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[14]_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.inst_addr_o[14] ),
    .A2(\i_snitch.pc_d[14] ));
 sg13g2_and3_1 \i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B  (.X(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y_sg13g2_and3_1_B_X ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_o21ai_1_A2_Y ),
    .C(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ));
 sg13g2_a21o_1 \i_snitch.pc_d[15]_sg13g2_a21o_1_A2  (.A2(\i_snitch.pc_d[15] ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1 ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_B1 ),
    .X(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X ));
 sg13g2_nor4_1 \i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D  (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ),
    .C(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ),
    .D(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D_Y ));
 sg13g2_a22oi_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[15] ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2308),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1 ),
    .A(net1396));
 sg13g2_xnor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1 ),
    .B(net2527));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C  (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .C(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1_sg13g2_o21ai_1_Y  (.B1(net2527),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_B1 ),
    .A1(\i_snitch.inst_addr_o[15] ),
    .A2(\i_snitch.inst_addr_o[16] ));
 sg13g2_a21oi_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1 ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand2_1_A_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1 ),
    .C(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2 ),
    .A(\i_snitch.inst_addr_o[15] ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ));
 sg13g2_nand3_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B ),
    .C(net64),
    .A(net2519),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nand3_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B ),
    .C(net63),
    .A(net2761),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A2(net2626));
 sg13g2_a21oi_2 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(net2852),
    .A1(net3019));
 sg13g2_or3_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X  (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B ),
    .C(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ),
    .X(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A_sg13g2_o21ai_1_Y  (.B1(net2528),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_B_sg13g2_inv_1_Y_A ),
    .A1(\i_snitch.inst_addr_o[13] ),
    .A2(\i_snitch.inst_addr_o[14] ));
 sg13g2_nor3_2 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ));
 sg13g2_nor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y  (.A(net2308),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2717),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2706),
    .C1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2613),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_xor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(net85),
    .X(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_and2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_B_X ),
    .X(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A_X ));
 sg13g2_xor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .X(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(net69));
 sg13g2_nor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B  (.A(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(net69),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2572),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .B1(net2538));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2586),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2593),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B  (.A(net2596),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2557),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2557),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2590),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2586),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ),
    .A(net2546),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_2 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .B(net2581),
    .A_N(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A(net2551),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X  (.A0(net2684),
    .A1(net2746),
    .S(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[16]_sg13g2_a221oi_1_A2  (.B2(\i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_B2 ),
    .C1(\i_snitch.pc_d[12]_sg13g2_mux2_1_A1_X ),
    .B1(\i_snitch.pc_d[22] ),
    .A1(\i_snitch.pc_d[16] ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_1 \i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_B2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_B2 ),
    .A(net1406));
 sg13g2_a22oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[16] ),
    .B1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2308),
    .A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1 ),
    .A(net1395));
 sg13g2_xnor2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1 ),
    .B(net2527));
 sg13g2_nand3_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1 ),
    .C(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2 ),
    .A(\i_snitch.inst_addr_o[16] ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2519),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_and3_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A ),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ),
    .C(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A ),
    .A(\i_snitch.inst_addr_o[15] ),
    .B(net2527));
 sg13g2_o21ai_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1  (.B1(net2762),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2 ),
    .B2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y ),
    .A2(net2629),
    .A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2_sg13g2_a21oi_1_Y  (.A1(net2991),
    .A2(net2852),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_B2 ),
    .B1(net2629));
 sg13g2_a21oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_and3_1_X_A ),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y  (.A(net2309),
    .B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2717),
    .B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2547),
    .C1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2613),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_inv_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ));
 sg13g2_nand2_2 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A ),
    .A(net2707),
    .B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .A2(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A(net2551),
    .B(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2749),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2715),
    .B(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2542),
    .Y(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2750),
    .A2(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[17] ),
    .A1(net2310),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2761),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2519));
 sg13g2_a221oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2  (.B2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .C1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ),
    .B1(net2761),
    .A1(net2965),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .A2(net2852));
 sg13g2_xnor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(net41));
 sg13g2_inv_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_A  (.Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_B1_sg13g2_a21oi_1_B1_A1 ),
    .A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[17] ),
    .B(net2528));
 sg13g2_nand2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_A1  (.A1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ),
    .B1(net2626));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2547),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_2 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.B1(net2538),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2572));
 sg13g2_o21ai_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2580),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2582),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2597),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .C1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2706),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2578));
 sg13g2_a21o_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .A1(net2580),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B_sg13g2_nor2_1_Y  (.A(net2592),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_or2_1_X_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A(net2584),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor2_1_B  (.A(net2584),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A1(net2594),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2562),
    .X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y  (.A1(net2600),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2600),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2594),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2581),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2577));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2598),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2596),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ),
    .A1(net2697),
    .B1(net2541),
    .X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2551),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(net2684),
    .A1(net2746),
    .S(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_and3_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_and3_1_C  (.X(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_B1 ),
    .A(\i_snitch.inst_addr_o[17] ),
    .B(net2313),
    .C(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor3_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[17] ),
    .B(net2306),
    .C(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A  (.A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ),
    .B(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_C_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_B1 ),
    .A(net893),
    .B(net2310));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2310),
    .Y(\i_snitch.pc_d[18] ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_xnor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1 ),
    .B(net2528));
 sg13g2_nor2b_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_B_N  (.A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B_N(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_A2 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2761),
    .C1(net2310),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2520),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2629),
    .A2(net2761),
    .A1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net2959),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_inv_4 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_inv_1_Y  (.A(net2853),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_nand3_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2 ),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_A_sg13g2_and4_1_C_B_sg13g2_nand4_1_D_Y ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand3_1_B_A ),
    .A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_a221oi_1_C1_A1_sg13g2_and4_1_X_A),
    .B(net3144));
 sg13g2_xnor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_or2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B ),
    .A(net75));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y  (.A1(net2577),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2580),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_or2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .B(net2599),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B_sg13g2_nor2_1_Y  (.A(net2592),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_B ));
 sg13g2_nor2_2 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2582),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2590),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2558),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2605),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2707),
    .A2(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2707),
    .B(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2604),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2558),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .A1(net2606),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2604),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2590),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2574),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A1(net2583),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B ),
    .Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2543),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A(net2697),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2553),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2749),
    .A2(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2614),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2 ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_Y ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nor3_1_A_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .A(net50),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_A  (.A(net50),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .X(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .B1(net2566));
 sg13g2_nor2b_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y  (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ),
    .B_N(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2573),
    .B1(net2538),
    .X(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2b_1 \i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_D_sg13g2_o21ai_1_Y_B1 ),
    .B(net2707),
    .A_N(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[18]_sg13g2_mux2_1_A1  (.A0(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[18] ),
    .S(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_A1 ),
    .X(\i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X ));
 sg13g2_a221oi_1 \i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1  (.B2(\i_snitch.inst_addr_o[27] ),
    .C1(\i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X ),
    .B1(net56),
    .A1(\i_snitch.inst_addr_o[22] ),
    .Y(\i_snitch.pc_d[18]_sg13g2_mux2_1_A1_X_sg13g2_a221oi_1_C1_Y ),
    .A2(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_inv_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2306),
    .Y(\i_snitch.pc_d[19] ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1166));
 sg13g2_a221oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2760),
    .C1(net2306),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1 ),
    .A2(net2520));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2760),
    .B(net71));
 sg13g2_nand2_2 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_a21o_1_B1_X ),
    .A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y  (.A(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_B_sg13g2_nor3_1_Y_B ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_a22oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2627),
    .A2(net2851),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ));
 sg13g2_nand4_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y  (.B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B ),
    .C(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C ),
    .A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .D(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D ));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_A ),
    .A(net2546),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(net2553),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_B_sg13g2_nand2_1_Y_B ),
    .A1(net2715),
    .A2(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C ),
    .A1(net2541),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(net2697),
    .A1(net2749),
    .S(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_C_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2707),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2614));
 sg13g2_xor2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(net66),
    .X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nor3_2 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .C(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X_B_sg13g2_nor2_1_B_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y ));
 sg13g2_a221oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_a221oi_1_B1  (.B2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y ),
    .C1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A_Y ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ),
    .Y(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_B ),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand3b_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C  (.B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ),
    .C(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C_Y ),
    .A_N(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_nand2b_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nor2b_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A  (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .B_N(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nor2b_1_A_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .A1(net2566),
    .A2(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor4_1_C_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2570),
    .B(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[273]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_B2_Y ));
 sg13g2_nor3_2 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.i_snitch_regfile.mem[304]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .C(\i_snitch.i_snitch_regfile.mem[51]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_xor2_1_B_X ),
    .A1(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_A_sg13g2_xor2_1_X_B_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2b_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B_N(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2  (.A1(net2546),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y  (.A1(net2551),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[300]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_A2_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2716),
    .B(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2577),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2586),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2574),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A1(net2586),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1 ),
    .B(\i_snitch.inst_addr_o[19] ));
 sg13g2_nor3_1 \i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[19] ),
    .B(net2306),
    .C(net62),
    .Y(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[1] ),
    .A1(net2301),
    .A2(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2755),
    .Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .B(net2515));
 sg13g2_nor2_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_Y ),
    .A1(net2718),
    .A2(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_B1 ),
    .A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .B(net2628));
 sg13g2_or2_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .B(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ),
    .A2(net2535),
    .Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_or2_1_X_B ),
    .B1(\i_snitch.inst_addr_o[1] ));
 sg13g2_nand3_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C  (.B(net2312),
    .C(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.inst_addr_o[1] ),
    .Y(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_B1 ));
 sg13g2_or3_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C  (.A(\i_snitch.inst_addr_o[1] ),
    .B(net2301),
    .C(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2 ),
    .X(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ));
 sg13g2_and4_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A  (.A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ),
    .D(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B_Y ),
    .X(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_B1 ),
    .A(net669),
    .B(net2301));
 sg13g2_mux2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X  (.A0(net1394),
    .A1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1 ),
    .S(net2313),
    .X(\i_snitch.pc_d[20] ));
 sg13g2_o21ai_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2  (.B1(\i_snitch.inst_addr_o[20] ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2_Y ),
    .A1(net2305),
    .A2(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1 ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .A1(net2717),
    .A2(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y  (.A1(net3134),
    .A2(net2851),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .B1(net2629));
 sg13g2_o21ai_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(net2626));
 sg13g2_xnor2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[20] ),
    .B(net2525));
 sg13g2_nand2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2761),
    .B(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2706),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ),
    .B(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .C1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2546),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21o_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A1(net2696),
    .B1(net2541),
    .X(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2551),
    .A2(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .A1(net2746),
    .S(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .X(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[20]_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[20]_sg13g2_or2_1_B_X ),
    .B(\i_snitch.pc_d[20] ),
    .A(\i_snitch.inst_addr_o[20] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[20]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[20]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[20]_sg13g2_or2_1_B_X ),
    .B2(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_A2_Y ),
    .A2(net419),
    .A1(\i_snitch.inst_addr_o[28] ));
 sg13g2_and2_1 \i_snitch.pc_d[20]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[20]_sg13g2_or2_1_B_X_sg13g2_a22oi_1_B1_Y ),
    .B(\i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1_Y ),
    .X(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2308),
    .Y(\i_snitch.pc_d[21] ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1242));
 sg13g2_a221oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2762),
    .C1(net2307),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1 ),
    .A2(net2519));
 sg13g2_a22oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2630),
    .A2(net2760),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(net2941),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_A2 ));
 sg13g2_xor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_xnor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.inst_addr_o[21] ),
    .B(net2526));
 sg13g2_a21oi_2 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.B1(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(net41));
 sg13g2_nand3_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A ),
    .A(net2706),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2577));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A(net2587),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1 ),
    .S(net2590),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net88),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y  (.A1(net2604),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2713),
    .A2(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2713),
    .B(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2605),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2704),
    .A2(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2705),
    .B(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y  (.A1(net2606),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2704),
    .A2(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B(net2704),
    .A_N(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2606),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .S(net2560),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net2603),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(net2711),
    .A2(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2711),
    .B(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .S(net2607),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2581),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2578));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2598),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net88),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .A1(net2604),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2605),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2596),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2551),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A(net2716),
    .B(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2543),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2697),
    .A2(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2746),
    .B(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2546),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2614));
 sg13g2_xnor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_and3_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C  (.X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B ),
    .C(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_inv_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B ),
    .A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_C ));
 sg13g2_nand3_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C  (.B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_B ),
    .C(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .A1(net46),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_a21o_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1  (.A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1_A1 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ),
    .X(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_B2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_a21o_1_B1_A1 ),
    .A(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X  (.B(net39),
    .A(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_and2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2b_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y  (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .B_N(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_and2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .A2(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .B1(net2566));
 sg13g2_a21oi_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2573),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_B  (.A(\i_snitch.inst_addr_o[21] ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[21] ),
    .B(net2308),
    .C(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[22] ));
 sg13g2_inv_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .A1(net2717),
    .A2(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_B1 ),
    .B(net2629),
    .A_N(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1  (.A1(net3096),
    .A2(net2852),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.inst_addr_o[22] ),
    .B(net2525));
 sg13g2_o21ai_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.inst_addr_o[21] ),
    .B(net2526));
 sg13g2_nor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2309),
    .B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2717),
    .B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .A1(net2614),
    .B1(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[22]_sg13g2_and2_1_X_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_B ),
    .A(\i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_B2 ),
    .B(net2308));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2309),
    .Y(\i_snitch.pc_d[23] ),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1372));
 sg13g2_a221oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2761),
    .C1(net2309),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2519),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y ),
    .B1(net2762),
    .B2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A2(net2852),
    .A1(net3090));
 sg13g2_nand2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_B1 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_B2_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[23] ),
    .B(net2525));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A2(net230));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2526),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.inst_addr_o[21] ),
    .A2(\i_snitch.inst_addr_o[22] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2613));
 sg13g2_xnor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_nor3_2 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nor4_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A ),
    .B(net39),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C ),
    .D(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y  (.B2(net2548),
    .C1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor2_2 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_a21oi_1_Y_B1 ),
    .B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_nand2b_1_Y_A_N ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_a221oi_1_Y_A1 ));
 sg13g2_nor4_2 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y ),
    .D(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1  (.B2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_B2 ),
    .C1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_A_Y ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_A1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_Y ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A ));
 sg13g2_nor3_2 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nor4_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A ),
    .B(net39),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C ),
    .D(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y  (.A(net2565),
    .B(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_Y  (.A(net2565),
    .B(net2548),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_C ));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_D ),
    .A(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_o21ai_1_A1  (.B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_C1_A1 ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_C ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_A ));
 sg13g2_nor3_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_nor3_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_X_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_A ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1 ),
    .B1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .X(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21o_1_X_A1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor3_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y  (.A(net2565),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_B1_A1 ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_inv_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C ),
    .A(net2548));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2569),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_A2  (.A1(net2569),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_A ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C ));
 sg13g2_nand4_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_Y  (.B(\i_snitch.i_snitch_regfile.mem[308]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[405]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .D(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nor3_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .A(net2547),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2573),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(net2539));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2589),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_A2  (.A1(net2584),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2579));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2599),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2594),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .S(net2554),
    .X(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2570),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand3_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_Y  (.B(net2554),
    .C(net2602),
    .A(net2599),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor4_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y  (.A(net2613),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B ),
    .C(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C ),
    .D(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2543),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2696),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2745),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2552),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D_sg13g2_nor2_1_Y  (.A(net75),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_nor4_1_Y_D ));
 sg13g2_o21ai_1 \i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X ));
 sg13g2_mux2_1 \i_snitch.pc_d[23]_sg13g2_mux2_1_A1  (.A0(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[23] ),
    .S(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_A1 ),
    .X(\i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1  (.A1(\i_snitch.inst_addr_o[24] ),
    .A2(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[23]_sg13g2_mux2_1_A1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2307),
    .Y(\i_snitch.pc_d[24] ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1346));
 sg13g2_a221oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2759),
    .C1(net2307),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2520),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2  (.B2(net2759),
    .C1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .A2(net2851));
 sg13g2_xor2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.inst_addr_o[24] ),
    .B(net2525));
 sg13g2_a21oi_2 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_or2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .B(net2526),
    .A(\i_snitch.inst_addr_o[23] ));
 sg13g2_a221oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1  (.B2(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ),
    .C1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_A_Y ),
    .A1(\i_snitch.inst_addr_o[24] ),
    .Y(\i_snitch.inst_addr_o[18]_sg13g2_a21o_1_A1_X_sg13g2_nand2_1_A_Y_sg13g2_a21oi_1_A1_Y_sg13g2_nand2b_1_A_N_B ),
    .A2(net2525));
 sg13g2_and2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.inst_addr_o[23] ),
    .B(net2526),
    .X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ));
 sg13g2_and2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ));
 sg13g2_a221oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .C1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2705),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21o_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(net2552),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .A1(net2745),
    .A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2543),
    .A2(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_A_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .B(net2696),
    .A_N(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a22oi_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2547),
    .A2(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2613));
 sg13g2_xnor2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21o_2 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ),
    .A1(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_nor2_1_A  (.A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ),
    .B(net2626),
    .Y(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_C1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[30] ),
    .B2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[24] ),
    .A1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_and2_1 \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y ),
    .B(\i_snitch.pc_d[28]_sg13g2_a22oi_1_A2_Y ),
    .X(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X ));
 sg13g2_nand4_1 \i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_A ),
    .C(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B ),
    .Y(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C_Y ),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2305),
    .Y(\i_snitch.pc_d[25] ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1197));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2  (.A1(\i_snitch.inst_addr_o[25] ),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2759),
    .C1(net2304),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2517),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2627),
    .A2(net2757),
    .A1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ),
    .B(net2853));
 sg13g2_xnor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[25] ),
    .B(net2523));
 sg13g2_a21o_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .A1(net41),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_and3_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ),
    .C(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2545),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2538));
 sg13g2_nand2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_A ),
    .A(net2703),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ),
    .A1(net75),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ));
 sg13g2_nor3_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y  (.A(net2611),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2542),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2696),
    .A2(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2745),
    .B(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2550),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(net2610),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_or3_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A  (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .C(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A_X ));
 sg13g2_xor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_nor2b_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_nor2b_1_B_N  (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .B_N(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor4_2 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nor3_1_Y_B_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D ),
    .C(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .D(net39));
 sg13g2_a21oi_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2548),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_and2_1_B_X ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_C ),
    .B1(net2565));
 sg13g2_and2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D_sg13g2_and2_1_X  (.A(net2569),
    .B(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nor4_1_Y_D ));
 sg13g2_o21ai_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_2 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_C_X ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.i_snitch_regfile.mem[408]_sg13g2_mux4_1_A0_X_sg13g2_a22oi_1_B1_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21o_1_B1_X ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[25] ),
    .B(net2305),
    .C(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2303),
    .Y(\i_snitch.pc_d[26] ),
    .B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1373));
 sg13g2_a221oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2757),
    .C1(net2303),
    .B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2517),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2757),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_or2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[26] ),
    .B(net2524));
 sg13g2_o21ai_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net41),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_A2 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21o_1_X_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.inst_addr_o[25] ),
    .B(net2523));
 sg13g2_a22oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2630),
    .A2(net2853),
    .A1(net3086));
 sg13g2_nand2_2 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2703),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2615));
 sg13g2_xor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_xor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .B(net103),
    .A_N(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N ));
 sg13g2_a221oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1 ),
    .C1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_and2_1_X_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_A2  (.A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A1 ),
    .B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1 ),
    .X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2545),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2695),
    .A2(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(net2540));
 sg13g2_a21o_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(net2550),
    .B1(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(net2749),
    .A2(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2684),
    .B(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a22oi_1 \i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1 ),
    .B2(\i_snitch.inst_addr_o[29] ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.inst_addr_o[26] ));
 sg13g2_nand2_1 \i_snitch.pc_d[26]_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[26]_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.pc_d[26] ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2303),
    .Y(\i_snitch.pc_d[27] ),
    .B1(net57));
 sg13g2_inv_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1075));
 sg13g2_a221oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2757),
    .C1(net2303),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1 ),
    .A2(net2517));
 sg13g2_nand2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2757),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2b_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A_N(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2523),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.inst_addr_o[25] ),
    .A2(\i_snitch.inst_addr_o[26] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2627),
    .A2(net2853),
    .A1(net3084));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2611));
 sg13g2_xor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A_Y ),
    .B2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N_Y ),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_a22oi_1_A1_A2 ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_nand2b_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A_N(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ));
 sg13g2_nand2b_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand3b_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y  (.B(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .C(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .A_N(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2_1_Y  (.A(net2564),
    .B(\i_snitch.i_snitch_regfile.mem[281]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_A_N ));
 sg13g2_inv_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_nor2_1_Y  (.A(net2568),
    .B(\i_snitch.i_snitch_regfile.mem[58]_sg13g2_a221oi_1_A1_Y_sg13g2_or3_1_C_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_nand3b_1_Y_B_sg13g2_inv_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2  (.B1(net2570),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A2(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_nand2b_1_B_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A_N(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y  (.A(net2611),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2716),
    .A2(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1  (.A2(net86),
    .A1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_B1  (.A1(net2716),
    .A2(net47),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A(net2549));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1 ),
    .A(net2748),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2698),
    .A2(\i_snitch.i_snitch_regfile.mem[283]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2540));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2545),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2699));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2578),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y  (.A(net2581),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2596),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(net2571),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y  (.A(net2592),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2554),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2562),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1 ),
    .X(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net2582),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2597),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1 ),
    .B2(net2579),
    .A2(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2544));
 sg13g2_o21ai_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1_sg13g2_o21ai_1_Y  (.B1(net2549),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a22oi_1_A2_B1 ),
    .A1(net2715),
    .A2(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ),
    .B1(net2539));
 sg13g2_a22oi_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .B1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2699),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C ),
    .A1(net2612));
 sg13g2_nor3_1 \i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[27] ),
    .B(net106),
    .C(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2304),
    .Y(\i_snitch.pc_d[28] ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1401));
 sg13g2_a221oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2758),
    .C1(net2304),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1 ),
    .A2(net2518));
 sg13g2_nand2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2758),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.inst_addr_o[28] ),
    .B(net2523));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(net72),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_or2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .B(net2523),
    .A(\i_snitch.inst_addr_o[27] ));
 sg13g2_and2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.inst_addr_o[27] ),
    .B(net2523),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2627),
    .A2(net2851),
    .A1(net3082));
 sg13g2_nand2_2 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2545),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2611));
 sg13g2_xor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_o21ai_1_Y_A2 ),
    .A2(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B1(net2539));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2588),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2595),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_or2_1_X_A ));
 sg13g2_mux2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2554),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .A(net2699),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2 ),
    .C1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2703),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2  (.A1(net2544),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1 ),
    .A1(net2610),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C ));
 sg13g2_a22oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2589),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2750),
    .A2(net2589));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2748),
    .A2(net2589),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B1(net2540));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2549),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2715),
    .A2(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2578),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2578),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2587),
    .A2(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .C1(net2585),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2591),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A1(net2559),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2560),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A(net88),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2554),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .B1(net2593));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net123),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2600),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .A1(net2716),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(net2550),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .A1(net2747),
    .A2(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_inv_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B2 ),
    .A(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2698),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .Y(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y_B ),
    .B1(net2540));
 sg13g2_a22oi_1 \i_snitch.pc_d[28]_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[28]_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1 ),
    .B2(\i_snitch.inst_addr_o[31] ),
    .A2(\i_snitch.pc_d[28] ),
    .A1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2303),
    .Y(\i_snitch.pc_d[29] ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1386));
 sg13g2_a221oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2757),
    .C1(net2304),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2517),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2627),
    .A2(net2758),
    .A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_A ),
    .A(net3080),
    .B(net2851));
 sg13g2_xnor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2b_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y  (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A ),
    .B_N(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_snitch.inst_addr_o[29] ),
    .B(net2524),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A ));
 sg13g2_a21oi_2 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_B_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2523),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.inst_addr_o[27] ),
    .A2(\i_snitch.inst_addr_o[28] ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2615),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand4_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A  (.B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .C(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y ),
    .D(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_or4_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D  (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_or3_1_A_X ),
    .B(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_C ),
    .D(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C ));
 sg13g2_nor2b_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y  (.A(net109),
    .B_N(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B  (.A(net109),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_and2_1_B_X ));
 sg13g2_nor3_2 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor3_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(net3144),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_B1_sg13g2_nor2b_1_Y_B_N ));
 sg13g2_or4_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D  (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_C ),
    .D(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X ));
 sg13g2_nand2_2 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_A ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ));
 sg13g2_nand3_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B_sg13g2_nand3_1_Y  (.B(net2923),
    .C(net2926),
    .A(net3033),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_B ));
 sg13g2_nand4_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D  (.B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_B ),
    .C(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1_Y ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y ),
    .D(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X ));
 sg13g2_xor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_and2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_xor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ),
    .A1(net2568),
    .A2(\i_snitch.i_snitch_regfile.mem[412]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.A1(net58),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2703),
    .C1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2545),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_A2  (.A1(net2711),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .B1(net2612));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .B1(net2539));
 sg13g2_inv_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2572),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2586),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2584),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y  (.A1(net2594),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2562),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net123),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2701),
    .A2(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2700),
    .B(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2601),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y  (.A1(net2701),
    .A2(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2700),
    .B(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_and2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2554),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .A1(net2600),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2700),
    .A2(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2700),
    .B(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2581),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_B1 ),
    .A1(net2594),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y  (.B1(net2574),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .A1(net2581),
    .A2(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_or3_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X  (.A(net2611),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C ),
    .X(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B ),
    .B1(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A(net2748),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y  (.A1(net2550),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C ),
    .B1(\i_snitch.i_snitch_regfile.mem[445]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A2 ),
    .A(net2716),
    .B(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[29]_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.pc_d[29] ));
 sg13g2_nand4_1 \i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A  (.B(\i_snitch.pc_d[26]_sg13g2_nand2_1_B_Y ),
    .C(\i_snitch.pc_d[16]_sg13g2_a221oi_1_A2_Y ),
    .A(\i_snitch.pc_d[15]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_D_Y ),
    .Y(\i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A_Y ),
    .D(\i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X  (.A0(net1378),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1 ),
    .S(net2312),
    .X(\i_snitch.pc_d[2] ));
 sg13g2_nand3_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C  (.B(net2312),
    .C(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1 ),
    .A(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1 ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_4 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.A(net2518),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_inv_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .B1(net2628),
    .B2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ),
    .A1(net2755));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .A(net84),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1  (.A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2 ),
    .B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .X(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_nand3_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2_sg13g2_nand3_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .C(net2535),
    .A(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_A1_A2 ));
 sg13g2_and3_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(net2535),
    .B(net3071),
    .C(\i_snitch.inst_addr_o[1] ));
 sg13g2_nor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor4_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_nor4_1_Y  (.A(\i_req_arb.data_i[37] ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .D(net2533),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .A2(net2535),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2755),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2612));
 sg13g2_nand4_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D  (.B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B ),
    .C(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_Y ),
    .D(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_xor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ),
    .X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A ));
 sg13g2_nand2_2 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ),
    .A(net2612),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B ));
 sg13g2_and2_2 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_and2_1_B  (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y ),
    .X(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B_Y ),
    .A(net43),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_A_N ),
    .A1(net2750),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y  (.A1(net2748),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1 ),
    .B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2610),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_o21ai_1_A2_B1_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A ));
 sg13g2_or2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ));
 sg13g2_and2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[64]_sg13g2_a221oi_1_A1_Y_sg13g2_nor4_1_C_Y_sg13g2_a21oi_1_B1_Y ),
    .B(net2602),
    .X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ),
    .X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(net2589),
    .B(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_A ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_nand2b_1_B  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A_sg13g2_xor2_1_X_B ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A_N(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ));
 sg13g2_nor3_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y  (.A(net2554),
    .B(net2602),
    .C(net2564),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net2608),
    .A2(net2570),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .B1(net2561));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A(net47),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_or2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ),
    .A(net47));
 sg13g2_xnor2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ),
    .A(net2593),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2554),
    .A2(net2600),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ),
    .B1(net2564));
 sg13g2_and2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y  (.A1(net2593),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A ),
    .B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2747),
    .A2(net47));
 sg13g2_a21oi_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2542),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1 ),
    .B1(net47));
 sg13g2_nand2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_X_A_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(net2695),
    .B(net2599));
 sg13g2_nand2_1 \i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .A(net2544),
    .B(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[2]_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_A ),
    .B(\i_snitch.pc_d[2] ),
    .Y(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2307),
    .Y(\i_snitch.pc_d[30] ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1 ),
    .A(net1390));
 sg13g2_xnor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1 ),
    .B(net2524));
 sg13g2_nand3b_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B  (.B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .C(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B_Y ),
    .A_N(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2759),
    .C1(net2304),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2517),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .A(net2759),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor2b_1_Y_A ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(\i_snitch.inst_addr_o[29] ),
    .B(net2523));
 sg13g2_a21oi_2 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A2(net54),
    .A1(net2611));
 sg13g2_xnor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_a221oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_B1 ),
    .C1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_A1 ),
    .A(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(net104));
 sg13g2_nor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(net104),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_xor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X  (.B(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_a21oi_1_Y  (.A1(net2570),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A_sg13g2_inv_1_A  (.Y(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_A ));
 sg13g2_a221oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .C1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(net2545),
    .A1(net2703),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2585),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2575),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .B1(net2593));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2561),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2 ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(net47),
    .A1(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .S(net2709),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2600),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(net2583),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2594),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .B1(net2539));
 sg13g2_a221oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2  (.B2(net2544),
    .C1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1 ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A1(net2699),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1 ),
    .A1(net2610),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net2542),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A ),
    .B1(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2695),
    .A2(net2556),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2747),
    .B(net2556),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2549),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .B1(net2556));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_C1_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .B(net2716));
 sg13g2_inv_2 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ));
 sg13g2_nor2_2 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A  (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y ),
    .B(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .A(net2610),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A2(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_a21o_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A1(net2748),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(net2550),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .A2(net2715));
 sg13g2_o21ai_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2542),
    .Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2750),
    .A2(\i_snitch.i_snitch_regfile.mem[286]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B2(net2629),
    .A2(net2851),
    .A1(net3078));
 sg13g2_nand2_1 \i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.inst_addr_o[30] ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_A1 ),
    .A2(net2303),
    .Y(\i_snitch.pc_d[31] ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_A1 ),
    .A(net696));
 sg13g2_a221oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(net2757),
    .C1(net2303),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2517),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2  (.B2(net2757),
    .C1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A_X ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A1(net3074),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .A2(net2853));
 sg13g2_xnor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.inst_addr_o[31] ),
    .B(net2524));
 sg13g2_nand2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_nand3b_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_o21ai_1_Y  (.B1(net2524),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .A1(\i_snitch.inst_addr_o[29] ),
    .A2(\i_snitch.inst_addr_o[30] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2611));
 sg13g2_inv_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2 ),
    .A(net77));
 sg13g2_xnor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .B(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ));
 sg13g2_xor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X  (.B(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y ),
    .A(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_A ));
 sg13g2_a21oi_2 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2  (.B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nor2b_1_A_Y ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_A2_Y ),
    .A2(net53),
    .A1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_xnor2_1_A_Y_sg13g2_nand2b_1_B_Y ));
 sg13g2_a221oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .C1(net2612),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21o_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .A1(net2748),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2550),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .A2(net2715));
 sg13g2_inv_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ),
    .A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_o21ai_1_A2  (.B1(net2542),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .A1(net2750),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_a221oi_1_Y_B2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2 ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2545),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2699));
 sg13g2_a221oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2  (.B2(net2699),
    .C1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2544),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y ),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ),
    .B(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B ),
    .A_N(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_nand2b_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_nand2b_1_Y_B ),
    .B(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_B1_X ),
    .A_N(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_or2_1_X_B ));
 sg13g2_inv_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_B1 ),
    .A2(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_X_sg13g2_xor2_1_B_X_sg13g2_xor2_1_B_X ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_A2_Y_sg13g2_inv_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2571),
    .A2(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21o_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2584),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(net2575),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1 ),
    .A1(net2589),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_Y_B ),
    .A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2599),
    .X(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y  (.B2(net2561),
    .C1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .A2(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1_sg13g2_nor2_1_Y  (.A(net2561),
    .B(net2601),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2701),
    .A2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2700),
    .B(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2700),
    .A2(\i_snitch.i_snitch_regfile.mem[159]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_B1_Y ));
 sg13g2_nor2b_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y  (.A(net2539),
    .B_N(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_B ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N ),
    .B1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_2 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B  (.A(net2576),
    .B(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_nor2_1_B_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .B(net2627),
    .X(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_and2_1_A_X ));
 sg13g2_nor3_1 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C  (.A(\i_snitch.inst_addr_o[31] ),
    .B(net2303),
    .C(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ));
 sg13g2_nor3_2 \i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_C_Y ),
    .B(\i_snitch.pc_d[29]_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_A_Y ),
    .C(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_Y_sg13g2_nand4_1_C_Y ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X  (.A2(net2301),
    .A1(net1119),
    .B1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[3] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B_Y ),
    .B2(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .A2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 ));
 sg13g2_inv_2 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 ),
    .A(net1119));
 sg13g2_and2_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X  (.A(net2312),
    .B(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1 ));
 sg13g2_nor3_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C  (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_A1 ),
    .B(net2302),
    .C(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ),
    .A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .B1(net2628),
    .B2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y ),
    .A1(net2756));
 sg13g2_xnor2_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2 ),
    .A(net82),
    .B(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21oi_2 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1  (.B1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A1(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N ));
 sg13g2_nor2b_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y  (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .B_N(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N ),
    .Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_and3_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_A ),
    .A(\i_req_arb.data_i[38] ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .C(net2535));
 sg13g2_a21o_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N_sg13g2_a21o_1_X  (.A2(net2535),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .B1(\i_req_arb.data_i[38] ),
    .X(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nor2b_1_Y_B_N ));
 sg13g2_nand2_1 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2755),
    .B(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[4] ),
    .A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net1393),
    .A2(net2301),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A ),
    .B1(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 ),
    .A_N(\i_req_arb.data_i[39] ));
 sg13g2_nor3_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .B(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ),
    .C(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .B1(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2518),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2755));
 sg13g2_nand3_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A ),
    .A1(net2540),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2_sg13g2_nand3_1_Y_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .B1(net2628),
    .B2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_A2 ),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2755));
 sg13g2_xnor2_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .A1(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ));
 sg13g2_nand3_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .C(net2535),
    .A(\i_req_arb.data_i[39] ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ));
 sg13g2_and3_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_A ),
    .A(\i_req_arb.data_i[39] ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .C(net2535));
 sg13g2_a21oi_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .A2(net122),
    .Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nor2_1_Y_B ),
    .B1(\i_req_arb.data_i[39] ));
 sg13g2_a22oi_1 \i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1 ),
    .B2(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ),
    .A2(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A ),
    .A1(\i_req_arb.data_i[39] ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .B(\i_snitch.pc_d[5] ),
    .Y(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A  (.A(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.pc_d[2]_sg13g2_nor2_1_B_Y ),
    .C(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_Y ),
    .Y(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y ));
 sg13g2_nand4_1 \i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y_sg13g2_nand4_1_D  (.B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N_Y ),
    .C(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_nand2_1_B_Y ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B_X ),
    .Y(\i_snitch.pc_d[11]_sg13g2_a21o_1_A2_X_sg13g2_nor4_1_A_D ),
    .D(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_Y_sg13g2_nor3_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5] ),
    .A1(net2301),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2518),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2755));
 sg13g2_nand2_2 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2544),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2612));
 sg13g2_xnor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_inv_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_C ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_nand3_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nand3_1_C  (.B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ),
    .C(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_B ));
 sg13g2_xor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_a21o_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_a21o_1_A2  (.A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21o_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B ),
    .A1(net115),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nor2b_2 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A  (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .B_N(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_B_N ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor3_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y  (.A(net2576),
    .B(net2564),
    .C(net59),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_A ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_B_N ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_B ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2572),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2584),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2594),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_and2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_and2_1_B  (.A(net2591),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .X(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .S(net2560),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net89),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(net2712),
    .A2(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2712),
    .B(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .A1(net2711),
    .A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2711),
    .B(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_mux2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .S(net89),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .A1(net2712),
    .A2(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2712),
    .B(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y  (.A1(net2704),
    .A2(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2704),
    .B(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2584),
    .B(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2574),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2587));
 sg13g2_nand2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A(net2590),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2557),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2607),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2607),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2557),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2606),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2604),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2595),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2587));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2560),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2603),
    .A2(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2603),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2560),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .A1(net65),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a221oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .C1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2699),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2571),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .B1(net2539));
 sg13g2_a21o_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .A1(net2580),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y  (.A1(net2592),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2555),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .A2(net123),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net123),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2592),
    .B(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2542),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2750),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2549),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(net2684),
    .A1(net2747),
    .S(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_xnor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1 ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B_sg13g2_a21oi_1_Y  (.A1(net2576),
    .A2(net61),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_B1_sg13g2_xnor2_1_A_B ),
    .B1(net2564));
 sg13g2_a22oi_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .B1(net2628),
    .B2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2756));
 sg13g2_xnor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .B(net45));
 sg13g2_xnor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .A(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .A(net3087),
    .B(net122));
 sg13g2_nor2_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B  (.A(net2301),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net1235),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ));
 sg13g2_inv_4 \i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.A(net645),
    .Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ));
 sg13g2_mux2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X  (.A0(net1361),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1 ),
    .S(net2312),
    .X(\i_snitch.pc_d[6] ));
 sg13g2_a21o_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2 ),
    .A1(net2518),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y ),
    .A(net2758),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B ),
    .A2(net2626));
 sg13g2_xor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2 ));
 sg13g2_nor3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_B  (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2 ));
 sg13g2_or2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1  (.A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2_sg13g2_a21o_1_X  (.A2(net2536),
    .A1(net3086),
    .B1(\i_req_arb.data_i[41] ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_B1_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B_Y ));
 sg13g2_nor4_2 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B ),
    .D(net2533));
 sg13g2_inv_2 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ),
    .A(net3085));
 sg13g2_nand4_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A  (.B(net3087),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B ),
    .Y(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_Y_sg13g2_a21oi_1_A1_B1 ),
    .D(net120));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C ));
 sg13g2_nor3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C  (.A(net96),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_C ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y ));
 sg13g2_a21o_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1  (.A2(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_A ),
    .A1(net93),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand3_1_C  (.B(net119),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_B ),
    .Y(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nor4_2 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nor4_1_Y  (.A(net3083),
    .B(net3077),
    .C(net3079),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C ),
    .D(net3081));
 sg13g2_nand2b_2 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A ),
    .A_N(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_nand3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N_sg13g2_nand3_1_Y  (.B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ),
    .C(net2926),
    .A(net3036),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nand2b_1_Y_A_N ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(net45),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_xnor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A(\i_req_arb.data_i[40] ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[5]_sg13g2_nor2_1_B_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y  (.A(net2718),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(net2544),
    .C1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2611),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B ),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nor4_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C ),
    .D(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_Y ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_C ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ));
 sg13g2_xor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_nand3b_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N  (.B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1 ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .A_N(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ),
    .B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_A2_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A ),
    .A1(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .A2(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_xor2_1_X_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ));
 sg13g2_inv_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2577),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A1 ),
    .B(net2586),
    .A_N(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .B1(net2578));
 sg13g2_or2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B ),
    .A(net2590));
 sg13g2_mux2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1 ),
    .S(net2560),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0 ),
    .A1(net2607),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2712),
    .A2(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2712),
    .B(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2607),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A1(net2704),
    .A2(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2704),
    .B(\i_snitch.i_snitch_regfile.mem[407]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1 ),
    .A1(net2603),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2702),
    .A2(\i_snitch.i_snitch_regfile.mem[152]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2702),
    .B(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_B  (.Y(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2603),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2603),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A1(net2702),
    .A2(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2702),
    .B(\i_snitch.i_snitch_regfile.mem[153]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2593),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2587));
 sg13g2_mux2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net88),
    .X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(net2606),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2 ),
    .A1(net75),
    .A2(\i_snitch.i_snitch_regfile.mem[148]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_or2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.i_snitch_regfile.mem[395]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .A(net2705));
 sg13g2_or2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .A(net89));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B ),
    .A1(net2704),
    .A2(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2705),
    .B(\i_snitch.i_snitch_regfile.mem[149]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .A1(net2604),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2707),
    .A2(\i_snitch.i_snitch_regfile.mem[141]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2708),
    .B(\i_snitch.i_snitch_regfile.mem[114]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2605),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A1(net2712),
    .A2(\i_snitch.i_snitch_regfile.mem[108]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y_B1 ),
    .A(net2713),
    .B(\i_snitch.i_snitch_regfile.mem[147]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2585),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_A ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B ),
    .A1(net2540),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2 ),
    .A1(net2747),
    .A2(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2695),
    .B(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C ),
    .A(\i_snitch.i_snitch_regfile.mem[38]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B_sg13g2_o21ai_1_Y  (.B1(net2550),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_nand3_1_Y_C_sg13g2_nand2_1_Y_B ),
    .A1(net2715),
    .A2(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand3_1 \i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C  (.B(net2312),
    .C(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1 ),
    .A(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_nand3_1_C_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[6]_sg13g2_o21ai_1_A2  (.B1(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_B1 ),
    .Y(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_Y ),
    .A1(\i_snitch.pc_d[6]_sg13g2_o21ai_1_A2_A1 ),
    .A2(\i_snitch.pc_d[6] ));
 sg13g2_a21o_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X  (.A2(net2302),
    .A1(net1196),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[7] ));
 sg13g2_a21oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1 ),
    .B1(net2302));
 sg13g2_nand2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1 ),
    .A(net2756),
    .B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ),
    .B(net2628));
 sg13g2_nand2_2 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ));
 sg13g2_nand2_2 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B ),
    .A(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2699),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2612));
 sg13g2_xnor2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nand3b_1_A_N_C ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_a21oi_2 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.B1(net2538),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2572));
 sg13g2_a221oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .C1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2544),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .A1(net2573),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2574),
    .B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2587));
 sg13g2_a21oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2591),
    .A2(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2590),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1 ),
    .A(net2591),
    .B(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2597),
    .A2(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2587));
 sg13g2_a21o_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ),
    .A1(net2695),
    .B1(net2540),
    .X(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2549),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_req_arb.data_i[42]_sg13g2_a221oi_1_A1_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(net2684),
    .A1(net2747),
    .S(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand3_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y  (.B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .A(net2518),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nand3_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B  (.B(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ),
    .C(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .A(net2756),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y ));
 sg13g2_or3_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ),
    .C(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ),
    .X(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y  (.A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_Y_A1 ),
    .A2(net45),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ),
    .B1(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_C ),
    .A1(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ),
    .A2(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ));
 sg13g2_nor3_1 \i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C  (.A(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ),
    .B(net2302),
    .C(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1 ),
    .Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_C_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a21oi_1_A2  (.A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8] ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_B1 ));
 sg13g2_nand4_1 \i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C  (.B(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_B_Y ),
    .C(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y ),
    .A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a21oi_1_A2_Y_sg13g2_nand4_1_C_Y ),
    .D(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_A2_Y ));
 sg13g2_a22oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[8] ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2 ),
    .A2(net2305),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_inv_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_A1 ),
    .A(net1405));
 sg13g2_and2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1 ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2 ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_and2_1_A_X ));
 sg13g2_nand3b_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y  (.B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B ),
    .C(net2517),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1 ),
    .A_N(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N ));
 sg13g2_nor2b_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N ),
    .B_N(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A_Y ));
 sg13g2_nor3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1  (.A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_Y ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ));
 sg13g2_a21o_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2_sg13g2_a21o_1_X  (.A2(net100),
    .A1(net3082),
    .B1(\i_req_arb.data_i[43] ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B ),
    .A(net3084),
    .B(net2536));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ),
    .A(\i_req_arb.data_i[42]_sg13g2_inv_1_A_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B ));
 sg13g2_nor3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ),
    .C(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B ));
 sg13g2_nand2b_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C ),
    .A_N(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_nor2_1_Y_B_sg13g2_xnor2_1_B_Y ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A_sg13g2_a21oi_1_Y  (.A1(net3082),
    .A2(net100),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_A ),
    .B1(\i_req_arb.data_i[43] ));
 sg13g2_and3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B_sg13g2_and3_1_X  (.X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nor2_1_Y_B ),
    .A(\i_req_arb.data_i[43] ),
    .B(net3082),
    .C(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_B ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2760),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2305));
 sg13g2_a21o_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .A1(net2613),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_nor4_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C  (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2 ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .D(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y ));
 sg13g2_nand2b_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_D ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_nor4_1_A_Y ),
    .A_N(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nand4_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B  (.B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_Y ),
    .D(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_inv_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_A ),
    .A(net102),
    .B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_A2_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_nor4_1_C_Y_sg13g2_nand4_1_B_C ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2 ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B ));
 sg13g2_nor3_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1_sg13g2_a21oi_1_Y  (.A1(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[262]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1_sg13g2_nand3_1_Y  (.B(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_o21ai_1_A2_Y ),
    .C(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor4_1_D_Y_sg13g2_or3_1_C_X ),
    .A(\i_snitch.i_snitch_regfile.mem[391]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_or3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A_sg13g2_or3_1_A  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B ),
    .X(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_and2_1_X_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B ));
 sg13g2_nor4_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C ),
    .D(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_B_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A ),
    .A2(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B ),
    .A1(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ));
 sg13g2_and2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ),
    .B(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_C_sg13g2_xnor2_1_Y_B_sg13g2_xor2_1_X_B ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_A_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_Y_C_sg13g2_nor4_1_Y_B ),
    .A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2b_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1  (.A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1_A2 ),
    .Y(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A ));
 sg13g2_nand2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1 ),
    .A(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_and3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B  (.X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B ),
    .C(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_nor3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y  (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C ),
    .A(\i_snitch.i_snitch_regfile.mem[138]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_A_sg13g2_nor3_1_Y_C_sg13g2_xnor2_1_Y_B ));
 sg13g2_nand3_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C  (.B(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_X ),
    .C(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_A1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y ));
 sg13g2_a21oi_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1  (.B1(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor3_1_A_Y_sg13g2_nand3b_1_C_Y ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y_sg13g2_a21oi_1_A1_Y ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_and3_1_B_X_sg13g2_nand3_1_C_Y ),
    .A1(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_B1_Y ));
 sg13g2_inv_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A ),
    .A(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ));
 sg13g2_xnor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_B_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B_sg13g2_xnor2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_2 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .A(net2546));
 sg13g2_a22oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2577));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2580),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2595),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2562),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2601),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ));
 sg13g2_nand2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2601),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2562),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2595),
    .B(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_inv_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nand2b_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B(net2586),
    .A_N(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y  (.A1(net2581),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2 ),
    .B1(net2578));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2590),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2557),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2604),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2604),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2557),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1 ));
 sg13g2_and2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X  (.A(net2596),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y  (.A1(net2559),
    .A2(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_or2_1_X_B_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2557),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_and2_1_X_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y  (.B2(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .C1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(net2705),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1 ),
    .A2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2543),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_inv_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2  (.B1(net2569),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .A1(net33),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y  (.A1(net2552),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .A1(net2745),
    .S(\i_snitch.i_snitch_regfile.mem[136]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_C1_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1  (.Y(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y ),
    .B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2 ),
    .B2(net2627),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor2b_1_A_Y ),
    .A1(net2758));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9] ),
    .A1(net2304),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2517),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2758));
 sg13g2_nand2_2 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_a22oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2547),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ),
    .A1(net2613));
 sg13g2_xor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X  (.B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2 ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ));
 sg13g2_and2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X  (.A(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A ));
 sg13g2_or2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B_sg13g2_or2_1_B  (.X(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_B1_sg13g2_a21oi_1_A1_A2 ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .A(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ));
 sg13g2_xnor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .A(net38),
    .B(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ));
 sg13g2_inv_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_inv_1_A  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_A1 ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y  (.A(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2  (.A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_A1 ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_B_sg13g2_a21oi_1_A2_Y ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_nor2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2577),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2585),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2592),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net2555),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net123),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(net2709),
    .A2(\i_snitch.i_snitch_regfile.mem[155]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2709),
    .B(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .A1(net2709),
    .A2(\i_snitch.i_snitch_regfile.mem[284]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2709),
    .B(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_mux4_1_A1_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_nand2b_1_A_N_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .A1(net2600),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2709),
    .A2(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_mux4_1_A0_X_sg13g2_a221oi_1_A2_Y_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_B1_X ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2710),
    .B(\i_snitch.i_snitch_regfile.mem[154]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .A(net2603),
    .B(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1 ),
    .B2(net2555),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y  (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .B(net2555),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1 ));
 sg13g2_nor2_2 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B  (.A(net2576),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(net2601));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1 ),
    .S(net2600),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0 ),
    .A1(net2701),
    .A2(\i_snitch.i_snitch_regfile.mem[158]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .A(net2700),
    .B(\i_snitch.i_snitch_regfile.mem[257]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1_sg13g2_mux2_1_X  (.A0(\i_snitch.i_snitch_regfile.mem[157]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .A1(net47),
    .S(net2709),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_B1_sg13g2_mux2_1_X_A1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2589),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_B2_sg13g2_a22oi_1_Y_B1_sg13g2_nor2b_1_Y_B_N_sg13g2_a21oi_1_Y_B1 ),
    .A2(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2582),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2596),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .S(net2558),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_A0  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_A_sg13g2_or2_1_X_B_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .S(net88),
    .X(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_nand3_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B ));
 sg13g2_mux2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X  (.A0(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .S(net89),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0 ),
    .A1(net75),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_or2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1_sg13g2_or2_1_X  (.X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A0_sg13g2_o21ai_1_Y_B1 ),
    .B(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .A(net2708));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1 ),
    .A1(net2707),
    .A2(\i_snitch.i_snitch_regfile.mem[400]_sg13g2_mux4_1_A0_1_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y ));
 sg13g2_nand2b_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A0_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1 ),
    .B(net2708),
    .A_N(\i_snitch.i_snitch_regfile.mem[143]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y  (.A1(net89),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2 ),
    .A1(net2712),
    .A2(\i_snitch.i_snitch_regfile.mem[142]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2713),
    .B(\i_snitch.i_snitch_regfile.mem[145]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net89),
    .B(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .A(net2597),
    .B(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2574),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1 ),
    .A1(net2582),
    .A2(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y  (.A1(net2705),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2573),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ),
    .B1(net2538));
 sg13g2_inv_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a21oi_1_Y_A2 ),
    .A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_B1_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_B1_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B1 ));
 sg13g2_a221oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2  (.B2(net2705),
    .C1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2547),
    .Y(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a21o_1_X_B1 ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_inv_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1 ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A ));
 sg13g2_a221oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y  (.B2(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_B_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_Y_C ),
    .C1(net2613),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2 ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2 ),
    .A1(net2745),
    .A2(net2548));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1_sg13g2_a21oi_1_Y  (.A1(net2696),
    .A2(net2548),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_A2_sg13g2_o21ai_1_Y_B1 ),
    .B1(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net2552),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_A2_sg13g2_a221oi_1_A2_C1_sg13g2_inv_1_Y_A_sg13g2_a221oi_1_Y_B1 ),
    .A1(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y ),
    .A2(\i_snitch.i_snitch_regfile.mem[150]_sg13g2_mux4_1_A0_1_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1 ),
    .A1(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y  (.A1(net2696),
    .A2(net37),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_A2 ),
    .B1(net2541));
 sg13g2_a21o_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .A1(net2552),
    .B1(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1 ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y  (.A1(net2716),
    .A2(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2 ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_nor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y  (.A(net2745),
    .B(\i_snitch.i_snitch_regfile.mem[41]_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a22oi_1_B2_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_B_sg13g2_a21oi_1_Y_B1_sg13g2_o21ai_1_Y_B1_sg13g2_a21o_1_X_A2_sg13g2_a21oi_1_Y_B1 ));
 sg13g2_a22oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .B1(net2627),
    .B2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2 ),
    .A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A1(net2758));
 sg13g2_xnor2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1 ),
    .A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ));
 sg13g2_a21o_2 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X  (.A2(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_A2 ),
    .A1(net45),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ));
 sg13g2_o21ai_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y  (.B1(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_A_sg13g2_a21oi_1_A1_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1 ),
    .A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21o_1_X_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3b_1_Y_A_N_sg13g2_nor3_1_Y_C_sg13g2_nand2b_1_B_Y ));
 sg13g2_a21oi_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1  (.A1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A ),
    .A2(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_nor3_1_B_Y ),
    .Y(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_or3_1_X_C_sg13g2_nor3_1_Y_B ),
    .B1(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_nand2_2 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_B ),
    .A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_C_sg13g2_a21oi_1_Y_A1 ),
    .B(\i_req_arb.data_i[44]_sg13g2_a21o_1_B1_X ));
 sg13g2_nand3_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C  (.B(net2312),
    .C(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_req_arb.data_i[44] ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ));
 sg13g2_nor2b_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N  (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_nor3_1_C_Y ),
    .B_N(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y ),
    .Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand3_1_C_Y_sg13g2_nor2b_1_B_N_Y ));
 sg13g2_or3_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C  (.A(\i_req_arb.data_i[44] ),
    .B(net2301),
    .C(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ));
 sg13g2_and4_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B  (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_a22oi_1_A2_Y ),
    .B(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X ),
    .C(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_A_X ),
    .D(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_A2_Y ),
    .X(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_or3_1_C_X_sg13g2_and4_1_B_X ));
 sg13g2_nand2_1 \i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_B1 ),
    .A(net1074),
    .B(net2304));
 sg13g2_o21ai_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[10] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2506),
    .Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2795),
    .B(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2795),
    .B(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2506),
    .Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1 ),
    .A(net560),
    .B(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[11] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2507),
    .Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2879),
    .B(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2879),
    .B(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2507),
    .Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1 ),
    .A(net573),
    .B(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y  (.B1(net556),
    .Y(\i_snitch.sb_d[12] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2503),
    .Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net3039),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net3039),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2504),
    .Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1 ),
    .A(net555),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand3_1 \i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y  (.B(\i_snitch.gpr_waddr[6] ),
    .C(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y),
    .A(\i_snitch.gpr_waddr[7] ),
    .Y(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y  (.B1(net558),
    .Y(\i_snitch.sb_d[13] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2505),
    .Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2861),
    .B(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2861),
    .B(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2505),
    .Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1 ),
    .A(net557),
    .B(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand3_1 \i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y  (.B(\i_snitch.gpr_waddr[6] ),
    .C(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .A(\i_snitch.gpr_waddr[7] ),
    .Y(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y  (.B1(net711),
    .Y(\i_snitch.sb_d[14] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2503),
    .Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2b_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B  (.Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .A_N(net2739));
 sg13g2_nor2_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2739),
    .B(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2739),
    .B(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2503),
    .Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_o21ai_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y  (.B1(net710),
    .Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1 ),
    .A1(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A2(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D));
 sg13g2_nand2_1 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_snitch.gpr_waddr[5] ),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y));
 sg13g2_nor2_2 \i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1 ),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D),
    .Y(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y  (.B1(net491),
    .Y(\i_snitch.sb_d[15] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2505),
    .Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2855),
    .B(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2855),
    .B(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2505),
    .Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1 ),
    .A(net490),
    .B(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_or2_1 \i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_or2_1_X  (.X(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_D),
    .A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y));
 sg13g2_o21ai_1 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[1] ),
    .A1(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1 ),
    .A2(net2292));
 sg13g2_nand2_2 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1 ),
    .A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1 ),
    .B(net2506),
    .Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2b_2 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B  (.Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .A_N(net2767));
 sg13g2_nor2_2 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2764),
    .B(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_2 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B  (.A(net2767),
    .B(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1 ),
    .C(net2506),
    .Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2b_1 \i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_B1 ),
    .B(net695),
    .A_N(net2767));
 sg13g2_o21ai_1 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[2] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ));
 sg13g2_nor2_2 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2506),
    .Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2b_2 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B  (.Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .B(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .A_N(net2783));
 sg13g2_nor2_2 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2782),
    .B(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_2 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2783),
    .B(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2506),
    .Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2b_1 \i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_B1 ),
    .B(net668),
    .A_N(net2785));
 sg13g2_o21ai_1 \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[3] ),
    .A1(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ),
    .A2(net2293));
 sg13g2_nor3_2 \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A  (.A(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1 ),
    .B(net2867),
    .C(net2506),
    .Y(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y ));
 sg13g2_nand2b_1 \i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2b_1_Y  (.Y(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_B1 ),
    .B(net593),
    .A_N(net2869));
 sg13g2_o21ai_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y  (.B1(net489),
    .Y(\i_snitch.sb_d[4] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_nor2_1_Y  (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ));
 sg13g2_nor2_2 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2503),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2887),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2887),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2503),
    .Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1 ),
    .A(net488),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[5] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2503),
    .Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2771),
    .B(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_2 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2773),
    .B(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2503),
    .Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1 ),
    .A(net540),
    .B(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[6] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_1_Y ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2503),
    .Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2790),
    .B(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2790),
    .B(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2504),
    .Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1 ),
    .A(net596),
    .B(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[7] ),
    .A1(net2293),
    .A2(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2504),
    .Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2874),
    .B(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2874),
    .B(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2504),
    .Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1 ),
    .A(net544),
    .B(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_2 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X),
    .B(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y  (.B1(net532),
    .Y(\i_snitch.sb_d[8] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_A ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2507),
    .Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2892),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(net2892),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2507),
    .Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1 ),
    .A(net531),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_o21ai_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y  (.B1(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1 ),
    .Y(\i_snitch.sb_d[9] ),
    .A1(net2292),
    .A2(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2 ));
 sg13g2_nand2_2 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .A(\i_snitch.gpr_waddr[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A1_sg13g2_nor2_1_B_Y ),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nand2_1_Y_B ));
 sg13g2_nor2_2 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A  (.A(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .B(net2507),
    .Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B  (.A(net2778),
    .B(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ),
    .Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ));
 sg13g2_nor3_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B  (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X),
    .B(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2 ),
    .C(net2507),
    .Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1 ),
    .A(net570),
    .B(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ));
 sg13g2_nand2_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A  (.Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .A(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .B(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y ));
 sg13g2_nand2_1 \i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y  (.Y(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B ),
    .A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y),
    .B(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_Y_B ));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3255),
    .D(\i_snitch.sb_d[10] ),
    .Q(\i_snitch.sb_q[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.sb_d[11] ),
    .Q(\i_snitch.sb_q[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[12] ),
    .Q(\i_snitch.sb_q[12] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.sb_d[13] ),
    .Q(\i_snitch.sb_q[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[14] ),
    .Q(\i_snitch.sb_q[14] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[15] ),
    .Q(\i_snitch.sb_q[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[1] ),
    .Q(\i_snitch.sb_q[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[2] ),
    .Q(\i_snitch.sb_q[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3254),
    .D(\i_snitch.sb_d[3] ),
    .Q(\i_snitch.sb_q[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_snitch.sb_d[4] ),
    .Q(\i_snitch.sb_q[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_snitch.sb_d[5] ),
    .Q(\i_snitch.sb_q[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3250),
    .D(\i_snitch.sb_d[6] ),
    .Q(\i_snitch.sb_q[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3220),
    .D(\i_snitch.sb_d[7] ),
    .Q(\i_snitch.sb_q[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 \i_snitch.sb_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.sb_d[8] ),
    .Q(\i_snitch.sb_q[8] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 \i_snitch.sb_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3223),
    .D(\i_snitch.sb_d[9] ),
    .Q(\i_snitch.sb_q[9] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.wake_up_q[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_mux2_1 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X  (.A0(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0 ),
    .A1(net1122),
    .S(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S ),
    .X(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_a21oi_1 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y  (.A1(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1 ),
    .A2(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ),
    .Y(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0 ),
    .B1(net1122));
 sg13g2_nor2_1 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2_sg13g2_nor2_1_Y  (.A(net553),
    .B(net545),
    .Y(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_A0_sg13g2_a21oi_1_Y_A2 ));
 sg13g2_mux2_1 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X  (.A0(net3),
    .A1(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1 ),
    .S(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ),
    .X(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S ));
 sg13g2_nand2_1 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y  (.Y(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1 ),
    .A(net3),
    .B(net645));
 sg13g2_dfrbpq_2 \i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(net646),
    .Q(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.wake_up_q[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_a22oi_1 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y  (.Y(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1 ),
    .B2(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2 ),
    .A2(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2 ),
    .A1(net553));
 sg13g2_or2_1 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X  (.X(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2 ),
    .B(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B ),
    .A(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ));
 sg13g2_nor3_1 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B_sg13g2_nor3_1_Y  (.A(net3),
    .B(net1122),
    .C(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ),
    .Y(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B ));
 sg13g2_nand2_1 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1_sg13g2_nand2_1_Y  (.Y(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B1 ),
    .A(net545),
    .B(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_A2_sg13g2_or2_1_X_B ));
 sg13g2_nor2_1 \i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y  (.A(net553),
    .B(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ),
    .Y(\i_snitch.wake_up_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a22oi_1_Y_B2 ));
 sg13g2_dfrbpq_2 \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\i_snitch.wake_up_q[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_nor3_1 \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y  (.A(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ),
    .B(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ),
    .C(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ),
    .Y(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_nor4_1 \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A_sg13g2_nor4_1_Y  (.A(net3),
    .B(net553),
    .C(net1122),
    .D(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X ),
    .Y(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_A ));
 sg13g2_and3_1 \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X  (.X(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B ),
    .A(net553),
    .B(net545),
    .C(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ));
 sg13g2_a21oi_1 \i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C_sg13g2_a21oi_1_Y  (.A1(net553),
    .A2(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_B_sg13g2_and3_1_X_C ),
    .Y(\i_snitch.wake_up_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor3_1_Y_C ),
    .B1(net545));
 sg13g2_nor4_1 \i_snitch.wake_up_q[2]_sg13g2_nor4_1_D  (.A(net3),
    .B(net553),
    .C(\i_snitch.wake_up_q[0] ),
    .D(net545),
    .Y(\i_snitch.wake_up_q[2]_sg13g2_nor4_1_D_Y ));
 sg13g2_nand2_1 \i_snitch.wake_up_q[2]_sg13g2_nor4_1_D_Y_sg13g2_nand2_1_B  (.Y(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q_D ),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X_sg13g2_nor3_1_B_Y_sg13g2_nand3_1_A_Y_sg13g2_nor4_1_A_Y_sg13g2_nand2_1_B_Y_sg13g2_or2_1_A_X_sg13g2_nand2_1_B_Y ),
    .B(\i_snitch.wake_up_q[2]_sg13g2_nor4_1_D_Y ));
 sg13g2_o21ai_1 req_data_valid_sg13g2_o21ai_1_Y (.B1(req_data_valid_sg13g2_o21ai_1_Y_B1),
    .Y(req_data_valid),
    .A1(net3053),
    .A2(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ));
 sg13g2_dfrbpq_2 \rsp_data_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(\rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_inv_1 \rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1354),
    .A2(net3064),
    .A1(net5));
 sg13g2_dfrbpq_2 \rsp_data_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3239),
    .D(\rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[10] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1336),
    .A2(net3066),
    .A1(net1322));
 sg13g2_dfrbpq_2 \rsp_data_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(\rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_inv_1 \rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1224));
 sg13g2_a22oi_1 \rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1223),
    .A2(net3064),
    .A1(\rsp_data_q[7] ));
 sg13g2_dfrbpq_2 \rsp_data_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(\rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[12] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_inv_1 \rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1306),
    .A2(net3065),
    .A1(net1183));
 sg13g2_dfrbpq_2 \rsp_data_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3239),
    .D(\rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[13] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1388),
    .A2(net3067),
    .A1(net1343));
 sg13g2_dfrbpq_2 \rsp_data_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(\rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[14] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1298));
 sg13g2_a22oi_1 \rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1297),
    .A2(net3066),
    .A1(\rsp_data_q[10] ));
 sg13g2_dfrbpq_2 \rsp_data_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3232),
    .D(\rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[15] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_inv_1 \rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1154));
 sg13g2_a22oi_1 \rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1153),
    .A2(net3064),
    .A1(\rsp_data_q[11] ));
 sg13g2_dfrbpq_2 \rsp_data_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(\rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[16] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_inv_1 \rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .A(net951));
 sg13g2_a22oi_1 \rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net950),
    .A2(net3063),
    .A1(\rsp_data_q[12] ));
 sg13g2_dfrbpq_2 \rsp_data_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[17] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_inv_1 \rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1350));
 sg13g2_a22oi_1 \rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1349),
    .A2(net3063),
    .A1(\rsp_data_q[13] ));
 sg13g2_dfrbpq_2 \rsp_data_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[18] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_inv_1 \rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1227));
 sg13g2_a22oi_1 \rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1226),
    .A2(net3067),
    .A1(\rsp_data_q[14] ));
 sg13g2_dfrbpq_2 \rsp_data_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3232),
    .D(\rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[19] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_inv_1 \rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1362),
    .A2(net3064),
    .A1(net1153));
 sg13g2_dfrbpq_2 \rsp_data_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3239),
    .D(\rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1382),
    .A2(net3064),
    .A1(net6));
 sg13g2_dfrbpq_2 \rsp_data_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[20] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_inv_1 \rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .A(net908));
 sg13g2_a22oi_1 \rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net907),
    .A2(net3063),
    .A1(\rsp_data_q[16] ));
 sg13g2_dfrbpq_2 \rsp_data_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3232),
    .D(\rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[21] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_inv_1 \rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1384),
    .A2(net3063),
    .A1(net1349));
 sg13g2_dfrbpq_2 \rsp_data_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3231),
    .D(\rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[22] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_inv_1 \rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1170));
 sg13g2_a22oi_1 \rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1169),
    .A2(net3063),
    .A1(\rsp_data_q[18] ));
 sg13g2_dfrbpq_2 \rsp_data_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[23] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_inv_1 \rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1272));
 sg13g2_a22oi_1 \rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1271),
    .A2(net3063),
    .A1(\rsp_data_q[19] ));
 sg13g2_dfrbpq_2 \rsp_data_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(\rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[24] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_inv_1 \rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1167),
    .A2(net3063),
    .A1(net907));
 sg13g2_dfrbpq_2 \rsp_data_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(\rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[25] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_inv_1 \rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1348));
 sg13g2_a22oi_1 \rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3062),
    .B2(net1347),
    .A2(net3063),
    .A1(\rsp_data_q[21] ));
 sg13g2_dfrbpq_2 \rsp_data_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3234),
    .D(\rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[26] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_inv_1 \rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3058),
    .B2(net1330),
    .A2(net3067),
    .A1(net1169));
 sg13g2_dfrbpq_2 \rsp_data_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3238),
    .D(\rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[27] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_inv_1 \rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3062),
    .B2(net1345),
    .A2(net3065),
    .A1(net1271));
 sg13g2_dfrbpq_2 \rsp_data_q[28]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3243),
    .D(\rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[28] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_inv_1 \rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1052));
 sg13g2_a22oi_1 \rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1051),
    .A2(net3065),
    .A1(\rsp_data_q[24] ));
 sg13g2_dfrbpq_2 \rsp_data_q[29]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(\rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[29] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_inv_1 \rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1294));
 sg13g2_a22oi_1 \rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1293),
    .A2(net3065),
    .A1(\rsp_data_q[25] ));
 sg13g2_dfrbpq_2 \rsp_data_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_inv_1 \rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1369),
    .A2(net3066),
    .A1(net7));
 sg13g2_dfrbpq_2 \rsp_data_q[30]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3244),
    .D(\rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[30] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_inv_1 \rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1158));
 sg13g2_a22oi_1 \rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1157),
    .A2(net3065),
    .A1(\rsp_data_q[26] ));
 sg13g2_dfrbpq_2 \rsp_data_q[31]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3239),
    .D(\rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[31] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1108));
 sg13g2_a22oi_1 \rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1107),
    .A2(net3065),
    .A1(\rsp_data_q[27] ));
 sg13g2_dfrbpq_2 \rsp_data_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_inv_1 \rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .A(\rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ));
 sg13g2_a22oi_1 \rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1381),
    .A2(net3066),
    .A1(net8));
 sg13g2_dfrbpq_2 \rsp_data_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(\rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_inv_1 \rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1264));
 sg13g2_a22oi_1 \rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1263),
    .A2(net3066),
    .A1(\rsp_data_q[0] ));
 sg13g2_dfrbpq_2 \rsp_data_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3240),
    .D(\rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1366));
 sg13g2_a22oi_1 \rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1365),
    .A2(net3065),
    .A1(\rsp_data_q[1] ));
 sg13g2_dfrbpq_2 \rsp_data_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(\rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_inv_1 \rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1323));
 sg13g2_a22oi_1 \rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1322),
    .A2(net3066),
    .A1(\rsp_data_q[2] ));
 sg13g2_dfrbpq_2 \rsp_data_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3237),
    .D(\rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_inv_1 \rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1300));
 sg13g2_a22oi_1 \rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3059),
    .B2(net1299),
    .A2(net3066),
    .A1(\rsp_data_q[3] ));
 sg13g2_dfrbpq_2 \rsp_data_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3241),
    .D(\rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_inv_1 \rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1184));
 sg13g2_a22oi_1 \rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3060),
    .B2(net1183),
    .A2(net3066),
    .A1(\rsp_data_q[4] ));
 sg13g2_dfrbpq_2 \rsp_data_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3239),
    .D(\rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\rsp_data_q[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_inv_1 \rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y  (.Y(\rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .A(net1344));
 sg13g2_a22oi_1 \rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y  (.Y(\rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .B1(net3061),
    .B2(net1343),
    .A2(net3065),
    .A1(\rsp_data_q[5] ));
 sg13g2_nor2b_1 rsp_data_ready_sg13g2_nor2b_1_Y (.A(net914),
    .B_N(net2),
    .Y(rsp_data_ready));
 sg13g2_and2_1 rsp_state_d_sg13g2_and2_1_X (.A(net4),
    .B(net3064),
    .X(rsp_state_d));
 sg13g2_dfrbpq_2 rsp_state_q_sg13g2_dfrbpq_1_Q (.RESET_B(net3232),
    .D(rsp_state_d),
    .Q(rsp_state_q),
    .CLK(clknet_leaf_36_clk));
 sg13g2_nor2_1 rsp_state_q_sg13g2_nor2_1_A (.A(net914),
    .B(net2),
    .Y(rsp_state_q_sg13g2_nor2_1_A_Y));
 sg13g2_a22oi_1 \shift_reg_q[0]_sg13g2_a22oi_1_A1  (.Y(uio_out_sg13g2_inv_1_Y_3_A),
    .B1(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_1_X ),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(\shift_reg_q[0] ));
 sg13g2_dfrbpq_1 \shift_reg_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3188),
    .D(net528),
    .Q(\shift_reg_q[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_a21oi_1 \shift_reg_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2732),
    .A2(\shift_reg_q[4]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[0]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[0]_sg13g2_nor2_1_A  (.A(net527),
    .B(net2732),
    .Y(\shift_reg_q[0]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[10]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[10]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(net468));
 sg13g2_dfrbpq_1 \shift_reg_q[10]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net469),
    .Q(\shift_reg_q[10] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[10]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2733),
    .A2(\shift_reg_q[14]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[10]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[10]_sg13g2_nor2_1_A  (.A(net468),
    .B(net2733),
    .Y(\shift_reg_q[10]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[11]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[11]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3055),
    .A2(net3045),
    .A1(\shift_reg_q[11] ));
 sg13g2_dfrbpq_1 \shift_reg_q[11]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net520),
    .Q(\shift_reg_q[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_a21oi_1 \shift_reg_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2731),
    .A2(\shift_reg_q[15]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[11]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[11]_sg13g2_nor2_1_A  (.A(net519),
    .B(net2731),
    .Y(\shift_reg_q[11]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[12]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[12]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3057),
    .A2(net3047),
    .A1(\shift_reg_q[12] ));
 sg13g2_dfrbpq_1 \shift_reg_q[12]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(net549),
    .Q(\shift_reg_q[12] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_a21oi_1 \shift_reg_q[12]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2735),
    .A2(\shift_reg_q[16]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[12]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[12]_sg13g2_nor2_1_A  (.A(net548),
    .B(net2735),
    .Y(\shift_reg_q[12]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[13]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[13]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3053),
    .A2(net3043),
    .A1(net476));
 sg13g2_dfrbpq_1 \shift_reg_q[13]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net477),
    .Q(\shift_reg_q[13] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_a21oi_1 \shift_reg_q[13]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2728),
    .A2(\shift_reg_q[17]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[13]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[13]_sg13g2_nor2_1_A  (.A(net476),
    .B(net2728),
    .Y(\shift_reg_q[13]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[14]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[14]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[14] ));
 sg13g2_dfrbpq_1 \shift_reg_q[14]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3198),
    .D(net487),
    .Q(\shift_reg_q[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2733),
    .A2(\shift_reg_q[18]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[14]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[14]_sg13g2_nor2_1_A  (.A(net486),
    .B(net2733),
    .Y(\shift_reg_q[14]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[15]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[15]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3055),
    .A2(net3045),
    .A1(net461));
 sg13g2_dfrbpq_1 \shift_reg_q[15]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3197),
    .D(net462),
    .Q(\shift_reg_q[15] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_a21oi_1 \shift_reg_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2731),
    .A2(\shift_reg_q[19]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[15]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[15]_sg13g2_nor2_1_A  (.A(net461),
    .B(net2732),
    .Y(\shift_reg_q[15]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[16]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[16]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3057),
    .A2(net3047),
    .A1(net546));
 sg13g2_dfrbpq_1 \shift_reg_q[16]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3230),
    .D(net547),
    .Q(\shift_reg_q[16] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_a21oi_1 \shift_reg_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2735),
    .A2(\shift_reg_q[20]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[16]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[16]_sg13g2_nor2_1_A  (.A(net546),
    .B(net2735),
    .Y(\shift_reg_q[16]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[17]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[17]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3053),
    .A2(net3043),
    .A1(\shift_reg_q[17] ));
 sg13g2_dfrbpq_1 \shift_reg_q[17]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net482),
    .Q(\shift_reg_q[17] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_a21oi_1 \shift_reg_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2729),
    .A2(\shift_reg_q[21]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[17]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[17]_sg13g2_nor2_1_A  (.A(net481),
    .B(net2729),
    .Y(\shift_reg_q[17]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[18]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[18]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[18] ));
 sg13g2_dfrbpq_1 \shift_reg_q[18]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net509),
    .Q(\shift_reg_q[18] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2733),
    .A2(\shift_reg_q[22]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[18]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[18]_sg13g2_nor2_1_A  (.A(net508),
    .B(net2734),
    .Y(\shift_reg_q[18]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[19]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[19]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3055),
    .A2(net3046),
    .A1(\shift_reg_q[19] ));
 sg13g2_dfrbpq_1 \shift_reg_q[19]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3197),
    .D(net499),
    .Q(\shift_reg_q[19] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_a21oi_1 \shift_reg_q[19]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2733),
    .A2(\shift_reg_q[23]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[19]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[19]_sg13g2_nor2_1_A  (.A(net498),
    .B(net2733),
    .Y(\shift_reg_q[19]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[1]_sg13g2_a22oi_1_A1  (.Y(uio_out_sg13g2_inv_1_Y_2_A),
    .B1(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(\shift_reg_q[1] ));
 sg13g2_dfrbpq_1 \shift_reg_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net536),
    .Q(\shift_reg_q[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_a21oi_1 \shift_reg_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2730),
    .A2(\shift_reg_q[5]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[1]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[1]_sg13g2_nor2_1_A  (.A(net535),
    .B(net2730),
    .Y(\shift_reg_q[1]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[20]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[20]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3057),
    .A2(net3047),
    .A1(net496));
 sg13g2_dfrbpq_1 \shift_reg_q[20]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3229),
    .D(net497),
    .Q(\shift_reg_q[20] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_a21oi_1 \shift_reg_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2735),
    .A2(\shift_reg_q[24]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[20]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[20]_sg13g2_nor2_1_A  (.A(net496),
    .B(net2736),
    .Y(\shift_reg_q[20]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[21]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[21]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3053),
    .A2(net3043),
    .A1(\shift_reg_q[21] ));
 sg13g2_dfrbpq_1 \shift_reg_q[21]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(net484),
    .Q(\shift_reg_q[21] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_a21oi_1 \shift_reg_q[21]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2728),
    .A2(\shift_reg_q[25]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[21]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[21]_sg13g2_nor2_1_A  (.A(net483),
    .B(net2728),
    .Y(\shift_reg_q[21]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[22]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[22]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[22] ));
 sg13g2_dfrbpq_1 \shift_reg_q[22]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3200),
    .D(net542),
    .Q(\shift_reg_q[22] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2734),
    .A2(\shift_reg_q[26]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[22]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[22]_sg13g2_nor2_1_A  (.A(net541),
    .B(net2734),
    .Y(\shift_reg_q[22]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[23]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[23]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[23] ));
 sg13g2_dfrbpq_1 \shift_reg_q[23]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net512),
    .Q(\shift_reg_q[23] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2734),
    .A2(\shift_reg_q[27]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[23]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[23]_sg13g2_nor2_1_A  (.A(net511),
    .B(net2734),
    .Y(\shift_reg_q[23]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[24]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[24]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3047),
    .A1(\shift_reg_q[24] ));
 sg13g2_dfrbpq_1 \shift_reg_q[24]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3229),
    .D(net530),
    .Q(\shift_reg_q[24] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_a21oi_1 \shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2735),
    .A2(\shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .Y(\shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[24]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .A1(net3172),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34] ));
 sg13g2_nor2_1 \shift_reg_q[24]_sg13g2_nor2_1_A  (.A(net529),
    .B(net2736),
    .Y(\shift_reg_q[24]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[25]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[25]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3053),
    .A2(net3044),
    .A1(\shift_reg_q[25] ));
 sg13g2_dfrbpq_1 \shift_reg_q[25]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3187),
    .D(net516),
    .Q(\shift_reg_q[25] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_a21oi_1 \shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2728),
    .A2(\shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .Y(\shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[25]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .A1(net3165),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35] ));
 sg13g2_nor2_1 \shift_reg_q[25]_sg13g2_nor2_1_A  (.A(net515),
    .B(net2728),
    .Y(\shift_reg_q[25]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[26]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[26]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[26] ));
 sg13g2_dfrbpq_1 \shift_reg_q[26]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3203),
    .D(net551),
    .Q(\shift_reg_q[26] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_a21oi_1 \shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2734),
    .A2(\shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .Y(\shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[26]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .A1(net3172),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36] ));
 sg13g2_nor2_1 \shift_reg_q[26]_sg13g2_nor2_1_A  (.A(net550),
    .B(net2734),
    .Y(\shift_reg_q[26]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[27]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[27]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3056),
    .A2(net3046),
    .A1(\shift_reg_q[27] ));
 sg13g2_dfrbpq_1 \shift_reg_q[27]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3199),
    .D(net615),
    .Q(\shift_reg_q[27] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_a21oi_1 \shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2737),
    .A2(\shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .Y(\shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[27]_sg13g2_nor2_1_A_Y ));
 sg13g2_o21ai_1 \shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y  (.B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_inv_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .Y(\shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_A2 ),
    .A1(net3170),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37] ));
 sg13g2_nor2_1 \shift_reg_q[27]_sg13g2_nor2_1_A  (.A(net614),
    .B(net2737),
    .Y(\shift_reg_q[27]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[2]_sg13g2_a22oi_1_A1  (.Y(uio_out_sg13g2_inv_1_Y_1_A),
    .B1(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(\shift_reg_q[2] ));
 sg13g2_dfrbpq_1 \shift_reg_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net480),
    .Q(\shift_reg_q[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_a21oi_1 \shift_reg_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2731),
    .A2(\shift_reg_q[6]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[2]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[2]_sg13g2_nor2_1_A  (.A(net479),
    .B(net2731),
    .Y(\shift_reg_q[2]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[3]_sg13g2_a22oi_1_A1  (.Y(uio_out_sg13g2_inv_1_Y_A),
    .B1(\shift_reg_q[0]_sg13g2_a22oi_1_A1_B1 ),
    .B2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_mux2_1_A1_1_X ),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(\shift_reg_q[3] ));
 sg13g2_dfrbpq_1 \shift_reg_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3188),
    .D(net522),
    .Q(\shift_reg_q[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_a21oi_1 \shift_reg_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2732),
    .A2(\shift_reg_q[7]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[3]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[3]_sg13g2_nor2_1_A  (.A(net521),
    .B(net2732),
    .Y(\shift_reg_q[3]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[4]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[4]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3057),
    .A2(net3047),
    .A1(net465));
 sg13g2_dfrbpq_1 \shift_reg_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3227),
    .D(net466),
    .Q(\shift_reg_q[4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_a21oi_1 \shift_reg_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2736),
    .A2(\shift_reg_q[8]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[4]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[4]_sg13g2_nor2_1_A  (.A(net465),
    .B(net2736),
    .Y(\shift_reg_q[4]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[5]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[5]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3053),
    .A2(net3044),
    .A1(net474));
 sg13g2_dfrbpq_1 \shift_reg_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3186),
    .D(net475),
    .Q(\shift_reg_q[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_a21oi_1 \shift_reg_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2730),
    .A2(\shift_reg_q[9]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[5]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[5]_sg13g2_nor2_1_A  (.A(net474),
    .B(net2730),
    .Y(\shift_reg_q[5]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[6]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[6]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3055),
    .A2(net3045),
    .A1(\shift_reg_q[6] ));
 sg13g2_dfrbpq_1 \shift_reg_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3197),
    .D(net507),
    .Q(\shift_reg_q[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_a21oi_1 \shift_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2733),
    .A2(\shift_reg_q[10]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[6]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[6]_sg13g2_nor2_1_A  (.A(net506),
    .B(net2731),
    .Y(\shift_reg_q[6]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[7]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[7]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3055),
    .A2(net3045),
    .A1(net492));
 sg13g2_dfrbpq_1 \shift_reg_q[7]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3195),
    .D(net493),
    .Q(\shift_reg_q[7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_a21oi_1 \shift_reg_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2731),
    .A2(\shift_reg_q[11]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[7]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[7]_sg13g2_nor2_1_A  (.A(net492),
    .B(net2731),
    .Y(\shift_reg_q[7]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[8]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[8]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3057),
    .A2(net3047),
    .A1(\shift_reg_q[8] ));
 sg13g2_dfrbpq_1 \shift_reg_q[8]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3229),
    .D(net504),
    .Q(\shift_reg_q[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_a21oi_1 \shift_reg_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2735),
    .A2(\shift_reg_q[12]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[8]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[8]_sg13g2_nor2_1_A  (.A(net503),
    .B(net2735),
    .Y(\shift_reg_q[8]_sg13g2_nor2_1_A_Y ));
 sg13g2_a22oi_1 \shift_reg_q[9]_sg13g2_a22oi_1_A1  (.Y(\shift_reg_q[9]_sg13g2_a22oi_1_A1_Y ),
    .B1(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_mux2_1_A1_1_X ),
    .B2(net3054),
    .A2(net3044),
    .A1(\shift_reg_q[9] ));
 sg13g2_dfrbpq_1 \shift_reg_q[9]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net539),
    .Q(\shift_reg_q[9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_a21oi_1 \shift_reg_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2728),
    .A2(\shift_reg_q[13]_sg13g2_a22oi_1_A1_Y ),
    .Y(\shift_reg_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\shift_reg_q[9]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \shift_reg_q[9]_sg13g2_nor2_1_A  (.A(net538),
    .B(net2728),
    .Y(\shift_reg_q[9]_sg13g2_nor2_1_A_Y ));
 sg13g2_dfrbpq_2 state_sg13g2_dfrbpq_1_Q (.RESET_B(net3184),
    .D(state_sg13g2_dfrbpq_1_Q_D),
    .Q(state),
    .CLK(clknet_leaf_1_clk));
 sg13g2_a21oi_1 state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y (.A1(net3053),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_B1 ),
    .Y(state_sg13g2_dfrbpq_1_Q_D),
    .B1(state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1));
 sg13g2_a21oi_1 state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_B1 (.A1(net1),
    .A2(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ),
    .Y(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B),
    .B1(state_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y_B1));
 sg13g2_inv_2 state_sg13g2_inv_1_A (.Y(state_sg13g2_inv_1_A_Y),
    .A(state));
 sg13g2_inv_1 strb_out_sg13g2_inv_1_Y (.Y(strb_out),
    .A(strb_out_sg13g2_inv_1_Y_A));
 sg13g2_a22oi_1 \strb_reg_q[0]_sg13g2_a22oi_1_A1  (.Y(strb_out_sg13g2_inv_1_Y_A),
    .B1(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B1 ),
    .B2(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B2 ),
    .A2(\cnt_q[2]_sg13g2_a22oi_1_B2_A2 ),
    .A1(\strb_reg_q[0] ));
 sg13g2_nor2_1 \strb_reg_q[0]_sg13g2_a22oi_1_A1_B1_sg13g2_nor2_1_Y  (.A(\i_req_register.data_o[5]_sg13g2_inv_1_A_Y ),
    .B(req_data_valid_sg13g2_o21ai_1_Y_B1),
    .Y(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \strb_reg_q[0]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3184),
    .D(net502),
    .Q(\strb_reg_q[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_a21oi_1 \strb_reg_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2730),
    .A2(\strb_reg_q[1]_sg13g2_a21oi_1_A1_Y ),
    .Y(\strb_reg_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[0]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[0]_sg13g2_nor2_1_A  (.A(net501),
    .B(net2730),
    .Y(\strb_reg_q[0]_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \strb_reg_q[1]_sg13g2_a21oi_1_A1  (.A1(\strb_reg_q[1] ),
    .A2(net3044),
    .Y(\strb_reg_q[1]_sg13g2_a21oi_1_A1_Y ),
    .B1(\strb_reg_q[0]_sg13g2_a22oi_1_A1_B2 ));
 sg13g2_dfrbpq_1 \strb_reg_q[1]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3185),
    .D(net526),
    .Q(\strb_reg_q[1] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_a21oi_1 \strb_reg_q[1]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2727),
    .A2(\strb_reg_q[2]_sg13g2_a21oi_1_A1_Y ),
    .Y(\strb_reg_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[1]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[1]_sg13g2_nor2_1_A  (.A(net525),
    .B(net2727),
    .Y(\strb_reg_q[1]_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \strb_reg_q[2]_sg13g2_a21oi_1_A1  (.A1(net517),
    .A2(net3043),
    .Y(\strb_reg_q[2]_sg13g2_a21oi_1_A1_Y ),
    .B1(\strb_reg_q[2]_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \strb_reg_q[2]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3185),
    .D(net518),
    .Q(\strb_reg_q[2] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_a21oi_1 \strb_reg_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2727),
    .A2(\strb_reg_q[3]_sg13g2_a21oi_1_A1_Y ),
    .Y(\strb_reg_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[2]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[2]_sg13g2_nor2_1_A  (.A(net517),
    .B(net2727),
    .Y(\strb_reg_q[2]_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \strb_reg_q[3]_sg13g2_a21oi_1_A1  (.A1(net459),
    .A2(net3043),
    .Y(\strb_reg_q[3]_sg13g2_a21oi_1_A1_Y ),
    .B1(\strb_reg_q[2]_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \strb_reg_q[3]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net460),
    .Q(\strb_reg_q[3] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_a21oi_1 \strb_reg_q[3]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2729),
    .A2(\strb_reg_q[4]_sg13g2_a21oi_1_A1_Y ),
    .Y(\strb_reg_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[3]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[3]_sg13g2_nor2_1_A  (.A(net459),
    .B(net2727),
    .Y(\strb_reg_q[3]_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \strb_reg_q[4]_sg13g2_a21oi_1_A1  (.A1(\strb_reg_q[4] ),
    .A2(net3043),
    .Y(\strb_reg_q[4]_sg13g2_a21oi_1_A1_Y ),
    .B1(\strb_reg_q[4]_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \strb_reg_q[4]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net473),
    .Q(\strb_reg_q[4] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_a21oi_1 \strb_reg_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(net2729),
    .A2(\strb_reg_q[5]_sg13g2_a21oi_1_A1_Y ),
    .Y(\strb_reg_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[4]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[4]_sg13g2_nor2_1_A  (.A(net472),
    .B(net2727),
    .Y(\strb_reg_q[4]_sg13g2_nor2_1_A_Y ));
 sg13g2_a21oi_1 \strb_reg_q[5]_sg13g2_a21oi_1_A1  (.A1(\strb_reg_q[5] ),
    .A2(net3043),
    .Y(\strb_reg_q[5]_sg13g2_a21oi_1_A1_Y ),
    .B1(\strb_reg_q[4]_sg13g2_a21oi_1_A1_B1 ));
 sg13g2_dfrbpq_1 \strb_reg_q[5]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(net443),
    .Q(\strb_reg_q[5] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_a21oi_1 \strb_reg_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y  (.A1(\strb_reg_q[6]_sg13g2_nand2_1_A_Y ),
    .A2(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ),
    .Y(\strb_reg_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .B1(\strb_reg_q[5]_sg13g2_nor2_1_A_Y ));
 sg13g2_nor2_1 \strb_reg_q[5]_sg13g2_nor2_1_A  (.A(\strb_reg_q[5] ),
    .B(net2727),
    .Y(\strb_reg_q[5]_sg13g2_nor2_1_A_Y ));
 sg13g2_dfrbpq_1 \strb_reg_q[6]_sg13g2_dfrbpq_1_Q  (.RESET_B(net3189),
    .D(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .Q(\strb_reg_q[6] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_nor2_1 \strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y  (.A(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ),
    .B(\strb_reg_q[6]_sg13g2_nor2_1_A_Y ),
    .Y(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D ));
 sg13g2_and2_1 \strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X  (.A(net2727),
    .B(net534),
    .X(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A ));
 sg13g2_nand2_1 \strb_reg_q[6]_sg13g2_nand2_1_A  (.Y(\strb_reg_q[6]_sg13g2_nand2_1_A_Y ),
    .A(net442),
    .B(net3043));
 sg13g2_nor2_1 \strb_reg_q[6]_sg13g2_nor2_1_A  (.A(net442),
    .B(net2729),
    .Y(\strb_reg_q[6]_sg13g2_nor2_1_A_Y ));
 sg13g2_dfrbpq_2 target_sel_q_sg13g2_dfrbpq_1_Q (.RESET_B(net3184),
    .D(net1027),
    .Q(target_sel_q),
    .CLK(clknet_leaf_6_clk));
 sg13g2_a21oi_1 target_sel_q_sg13g2_dfrbpq_1_Q_D_sg13g2_a21oi_1_Y (.A1(target_sel_q_sg13g2_nor2_1_A_B),
    .A2(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_a21oi_1_A2_Y ),
    .Y(target_sel_q_sg13g2_dfrbpq_1_Q_D),
    .B1(target_sel_q_sg13g2_nor2_1_A_Y));
 sg13g2_nand2_1 target_sel_q_sg13g2_nand2_1_B (.Y(target_sel_q_sg13g2_nand2_1_B_Y),
    .A(net914),
    .B(net1026));
 sg13g2_nand2b_2 target_sel_q_sg13g2_nand2b_1_A_N (.Y(target_sel_q_sg13g2_nand2b_1_A_N_Y),
    .B(net914),
    .A_N(target_sel_q));
 sg13g2_nand2b_2 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N (.Y(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y),
    .B(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nand2_1_Y_B ),
    .A_N(target_sel_q_sg13g2_nand2b_1_A_N_Y));
 sg13g2_nor2_1 target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A (.A(target_sel_q_sg13g2_nand2b_1_A_N_Y),
    .B(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_B),
    .Y(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_Y));
 sg13g2_nor2_1 target_sel_q_sg13g2_nor2_1_A (.A(net1026),
    .B(target_sel_q_sg13g2_nor2_1_A_B),
    .Y(target_sel_q_sg13g2_nor2_1_A_Y));
 sg13g2_nor2_1 target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y (.A(req_data_valid_sg13g2_o21ai_1_Y_B1),
    .B(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B),
    .Y(target_sel_q_sg13g2_nor2_1_A_B));
 sg13g2_nand3b_1 target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B (.B(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B),
    .C(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .Y(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B_Y),
    .A_N(net3164));
 sg13g2_tiehi heichips25_snitch_wrapper_26 (.L_HI(net26));
 sg13g2_tiehi heichips25_snitch_wrapper_27 (.L_HI(net27));
 sg13g2_tiehi heichips25_snitch_wrapper_28 (.L_HI(net28));
 sg13g2_tiehi heichips25_snitch_wrapper_29 (.L_HI(net29));
 sg13g2_tiehi heichips25_snitch_wrapper_30 (.L_HI(net30));
 sg13g2_tiehi heichips25_snitch_wrapper_31 (.L_HI(net31));
 sg13g2_tiehi heichips25_snitch_wrapper_32 (.L_HI(net32));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 uio_out_sg13g2_buf_1_X (.A(\i_req_register.data_o[42] ),
    .X(net13));
 sg13g2_buf_1 uio_out_sg13g2_buf_1_X_1 (.A(\i_req_register.data_o[43] ),
    .X(net14));
 sg13g2_buf_1 uio_out_sg13g2_buf_1_X_2 (.A(\i_req_register.data_o[44] ),
    .X(net15));
 sg13g2_buf_1 uio_out_sg13g2_buf_1_X_3 (.A(\i_req_register.data_o[45] ),
    .X(net16));
 sg13g2_inv_1 uio_out_sg13g2_inv_1_Y (.Y(net12),
    .A(uio_out_sg13g2_inv_1_Y_A));
 sg13g2_inv_1 uio_out_sg13g2_inv_1_Y_1 (.Y(net11),
    .A(uio_out_sg13g2_inv_1_Y_1_A));
 sg13g2_inv_1 uio_out_sg13g2_inv_1_Y_2 (.Y(net10),
    .A(uio_out_sg13g2_inv_1_Y_2_A));
 sg13g2_inv_1 uio_out_sg13g2_inv_1_Y_3 (.Y(net9),
    .A(uio_out_sg13g2_inv_1_Y_3_A));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X (.A(req_data_valid),
    .X(net17));
 sg13g2_buf_8 uo_out_sg13g2_buf_1_X_1 (.A(net3064),
    .X(net18));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X_2 (.A(strb_out),
    .X(net19));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X_3 (.A(\i_req_register.data_o[5] ),
    .X(net20));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X_4 (.A(\i_req_register.data_o[38] ),
    .X(net21));
 sg13g2_buf_8 uo_out_sg13g2_buf_1_X_5 (.A(\i_req_register.data_o[39] ),
    .X(net22));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X_6 (.A(\i_req_register.data_o[40] ),
    .X(net23));
 sg13g2_buf_1 uo_out_sg13g2_buf_1_X_7 (.A(\i_req_register.data_o[41] ),
    .X(net24));
 sg13g2_buf_16 fanout2237 (.X(net2237),
    .A(net2238));
 sg13g2_buf_16 fanout2238 (.X(net2238),
    .A(net2241));
 sg13g2_buf_16 fanout2239 (.X(net2239),
    .A(net68));
 sg13g2_buf_16 fanout2240 (.X(net2240),
    .A(net68));
 sg13g2_buf_8 fanout2241 (.A(\i_snitch.pc_d[24]_sg13g2_a22oi_1_A2_Y_sg13g2_and2_1_A_X_sg13g2_nand4_1_C_Y ),
    .X(net2241));
 sg13g2_buf_8 fanout2242 (.A(net2243),
    .X(net2242));
 sg13g2_buf_8 fanout2243 (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .X(net2243));
 sg13g2_buf_8 fanout2244 (.A(net2245),
    .X(net2244));
 sg13g2_buf_8 fanout2245 (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2245));
 sg13g2_buf_8 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_8 fanout2247 (.A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2247));
 sg13g2_buf_8 fanout2248 (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y ),
    .X(net2248));
 sg13g2_buf_8 fanout2249 (.A(\i_snitch.pc_d[23]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_A1_Y ),
    .X(net2249));
 sg13g2_buf_8 fanout2250 (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .X(net2250));
 sg13g2_buf_8 fanout2251 (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .X(net2251));
 sg13g2_buf_8 fanout2252 (.A(net2253),
    .X(net2252));
 sg13g2_buf_8 fanout2253 (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2253));
 sg13g2_buf_8 fanout2254 (.A(net2255),
    .X(net2254));
 sg13g2_buf_8 fanout2255 (.A(\i_snitch.pc_d[26]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2255));
 sg13g2_buf_8 fanout2256 (.A(net2257),
    .X(net2256));
 sg13g2_buf_8 fanout2257 (.A(\i_snitch.pc_d[24]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .X(net2257));
 sg13g2_buf_8 fanout2258 (.A(net2259),
    .X(net2258));
 sg13g2_buf_8 fanout2259 (.A(\i_snitch.pc_d[22]_sg13g2_and2_1_X_A_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(net2259));
 sg13g2_buf_8 fanout2260 (.A(net2261),
    .X(net2260));
 sg13g2_buf_8 fanout2261 (.A(\i_snitch.pc_d[20]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2261));
 sg13g2_buf_8 fanout2262 (.A(net2263),
    .X(net2262));
 sg13g2_buf_8 fanout2263 (.A(\i_snitch.pc_d[16]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_o21ai_1_A1_Y_sg13g2_a22oi_1_B1_Y ),
    .X(net2263));
 sg13g2_buf_8 fanout2264 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .X(net2264));
 sg13g2_buf_8 fanout2265 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_B_sg13g2_nand3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_a21oi_1_B1_Y ),
    .X(net2265));
 sg13g2_buf_8 fanout2266 (.A(net2267),
    .X(net2266));
 sg13g2_buf_8 fanout2267 (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_nand2_1_B_Y ),
    .X(net2267));
 sg13g2_buf_8 fanout2268 (.A(net2269),
    .X(net2268));
 sg13g2_buf_8 fanout2269 (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2269));
 sg13g2_buf_8 fanout2270 (.A(net2271),
    .X(net2270));
 sg13g2_buf_8 fanout2271 (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2271));
 sg13g2_buf_8 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_8 fanout2273 (.A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_a22oi_1_A2_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2273));
 sg13g2_buf_8 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_8 fanout2275 (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_A_Y ),
    .X(net2275));
 sg13g2_buf_8 fanout2276 (.A(net2277),
    .X(net2276));
 sg13g2_buf_8 fanout2277 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_Y ),
    .X(net2277));
 sg13g2_buf_8 fanout2278 (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y ),
    .X(net2278));
 sg13g2_buf_8 fanout2279 (.A(\i_snitch.pc_d[8]_sg13g2_a22oi_1_Y_B2_sg13g2_a21oi_1_Y_A2_sg13g2_a22oi_1_B1_Y ),
    .X(net2279));
 sg13g2_buf_8 fanout2280 (.A(net2281),
    .X(net2280));
 sg13g2_buf_8 fanout2281 (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_nand3_1_C_Y_sg13g2_and2_1_B_X ),
    .X(net2281));
 sg13g2_buf_8 fanout2282 (.A(net2283),
    .X(net2282));
 sg13g2_buf_8 fanout2283 (.A(\i_snitch.pc_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2283));
 sg13g2_buf_8 fanout2284 (.A(net2285),
    .X(net2284));
 sg13g2_buf_8 fanout2285 (.A(\i_snitch.pc_d[7]_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y_sg13g2_nand2_1_A_Y ),
    .X(net2285));
 sg13g2_buf_8 fanout2286 (.A(net2287),
    .X(net2286));
 sg13g2_buf_8 fanout2287 (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_nand2_1_B_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2287));
 sg13g2_buf_8 fanout2288 (.A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .X(net2288));
 sg13g2_buf_8 fanout2289 (.A(\i_snitch.pc_d[17]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_a221oi_1_B2_Y ),
    .X(net2289));
 sg13g2_buf_8 fanout2290 (.A(net2291),
    .X(net2290));
 sg13g2_buf_8 fanout2291 (.A(\i_snitch.pc_d[13]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_o21ai_1_A2_Y ),
    .X(net2291));
 sg13g2_buf_8 fanout2292 (.A(net2293),
    .X(net2292));
 sg13g2_buf_8 fanout2293 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_Y_sg13g2_nand3_1_C_Y ),
    .X(net2293));
 sg13g2_buf_8 fanout2294 (.A(net2295),
    .X(net2294));
 sg13g2_buf_8 fanout2295 (.A(net2298),
    .X(net2295));
 sg13g2_buf_8 fanout2296 (.A(net2297),
    .X(net2296));
 sg13g2_buf_8 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_8 fanout2298 (.A(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2_1_A_Y),
    .X(net2298));
 sg13g2_buf_8 fanout2299 (.A(net2300),
    .X(net2299));
 sg13g2_buf_8 fanout2300 (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .X(net2300));
 sg13g2_buf_8 fanout2301 (.A(net2302),
    .X(net2301));
 sg13g2_buf_8 fanout2302 (.A(net2311),
    .X(net2302));
 sg13g2_buf_8 fanout2303 (.A(net2304),
    .X(net2303));
 sg13g2_buf_8 fanout2304 (.A(net106),
    .X(net2304));
 sg13g2_buf_8 fanout2305 (.A(net2307),
    .X(net2305));
 sg13g2_buf_1 fanout2306 (.A(net2307),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(net106),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(net2309),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(net2310),
    .X(net2309));
 sg13g2_buf_2 fanout2310 (.A(net106),
    .X(net2310));
 sg13g2_buf_8 fanout2311 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_or2_1_B_X ),
    .X(net2311));
 sg13g2_buf_8 fanout2312 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ),
    .X(net2312));
 sg13g2_buf_1 fanout2313 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y ),
    .X(net2313));
 sg13g2_buf_8 fanout2314 (.A(net2315),
    .X(net2314));
 sg13g2_buf_8 fanout2315 (.A(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2315));
 sg13g2_buf_8 fanout2316 (.A(net2320),
    .X(net2316));
 sg13g2_buf_8 fanout2317 (.A(net2319),
    .X(net2317));
 sg13g2_buf_8 fanout2318 (.A(net2319),
    .X(net2318));
 sg13g2_buf_8 fanout2319 (.A(net2320),
    .X(net2319));
 sg13g2_buf_8 fanout2320 (.A(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2320));
 sg13g2_buf_8 fanout2321 (.A(net2322),
    .X(net2321));
 sg13g2_buf_8 fanout2322 (.A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2322));
 sg13g2_buf_8 fanout2323 (.A(net2327),
    .X(net2323));
 sg13g2_buf_8 fanout2324 (.A(net2327),
    .X(net2324));
 sg13g2_buf_8 fanout2325 (.A(net2326),
    .X(net2325));
 sg13g2_buf_8 fanout2326 (.A(net2327),
    .X(net2326));
 sg13g2_buf_8 fanout2327 (.A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2327));
 sg13g2_buf_8 fanout2328 (.A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2328));
 sg13g2_buf_8 fanout2329 (.A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2329));
 sg13g2_buf_8 fanout2330 (.A(net2333),
    .X(net2330));
 sg13g2_buf_8 fanout2331 (.A(net2333),
    .X(net2331));
 sg13g2_buf_8 fanout2332 (.A(net2333),
    .X(net2332));
 sg13g2_buf_8 fanout2333 (.A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2333));
 sg13g2_buf_8 fanout2334 (.A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2334));
 sg13g2_buf_8 fanout2335 (.A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2335));
 sg13g2_buf_8 fanout2336 (.A(net2339),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(net2338),
    .X(net2337));
 sg13g2_buf_8 fanout2338 (.A(net2339),
    .X(net2338));
 sg13g2_buf_8 fanout2339 (.A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2339));
 sg13g2_buf_8 fanout2340 (.A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2341));
 sg13g2_buf_8 fanout2342 (.A(net2346),
    .X(net2342));
 sg13g2_buf_8 fanout2343 (.A(net2346),
    .X(net2343));
 sg13g2_buf_8 fanout2344 (.A(net2346),
    .X(net2344));
 sg13g2_buf_8 fanout2345 (.A(net2346),
    .X(net2345));
 sg13g2_buf_8 fanout2346 (.A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2346));
 sg13g2_buf_8 fanout2347 (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2347));
 sg13g2_buf_8 fanout2348 (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2348));
 sg13g2_buf_8 fanout2349 (.A(net2352),
    .X(net2349));
 sg13g2_buf_8 fanout2350 (.A(net2351),
    .X(net2350));
 sg13g2_buf_8 fanout2351 (.A(net2352),
    .X(net2351));
 sg13g2_buf_8 fanout2352 (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2352));
 sg13g2_buf_8 fanout2353 (.A(net2354),
    .X(net2353));
 sg13g2_buf_8 fanout2354 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2354));
 sg13g2_buf_8 fanout2355 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2355));
 sg13g2_buf_8 fanout2356 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2356));
 sg13g2_buf_8 fanout2357 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2357));
 sg13g2_buf_8 fanout2358 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2358));
 sg13g2_buf_8 fanout2359 (.A(net2360),
    .X(net2359));
 sg13g2_buf_8 fanout2360 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2360));
 sg13g2_buf_8 fanout2361 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2361));
 sg13g2_buf_8 fanout2362 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2362));
 sg13g2_buf_8 fanout2363 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2363));
 sg13g2_buf_2 fanout2364 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2364));
 sg13g2_buf_8 fanout2365 (.A(net2366),
    .X(net2365));
 sg13g2_buf_8 fanout2366 (.A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2366));
 sg13g2_buf_8 fanout2367 (.A(net2371),
    .X(net2367));
 sg13g2_buf_8 fanout2368 (.A(net2370),
    .X(net2368));
 sg13g2_buf_8 fanout2369 (.A(net2371),
    .X(net2369));
 sg13g2_buf_8 fanout2370 (.A(net2371),
    .X(net2370));
 sg13g2_buf_8 fanout2371 (.A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2371));
 sg13g2_buf_8 fanout2372 (.A(net2376),
    .X(net2372));
 sg13g2_buf_8 fanout2373 (.A(net2375),
    .X(net2373));
 sg13g2_buf_8 fanout2374 (.A(net2376),
    .X(net2374));
 sg13g2_buf_8 fanout2375 (.A(net2376),
    .X(net2375));
 sg13g2_buf_8 fanout2376 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2376));
 sg13g2_buf_8 fanout2377 (.A(net2378),
    .X(net2377));
 sg13g2_buf_8 fanout2378 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2378));
 sg13g2_buf_8 fanout2379 (.A(net2380),
    .X(net2379));
 sg13g2_buf_8 fanout2380 (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2380));
 sg13g2_buf_8 fanout2381 (.A(net2383),
    .X(net2381));
 sg13g2_buf_8 fanout2382 (.A(net2383),
    .X(net2382));
 sg13g2_buf_8 fanout2383 (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2383));
 sg13g2_buf_8 fanout2384 (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2384));
 sg13g2_buf_8 fanout2385 (.A(net2386),
    .X(net2385));
 sg13g2_buf_8 fanout2386 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2386));
 sg13g2_buf_8 fanout2387 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2387));
 sg13g2_buf_8 fanout2388 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2388));
 sg13g2_buf_8 fanout2389 (.A(net2391),
    .X(net2389));
 sg13g2_buf_8 fanout2390 (.A(net2391),
    .X(net2390));
 sg13g2_buf_8 fanout2391 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2391));
 sg13g2_buf_8 fanout2392 (.A(net2393),
    .X(net2392));
 sg13g2_buf_8 fanout2393 (.A(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2393));
 sg13g2_buf_8 fanout2394 (.A(net2398),
    .X(net2394));
 sg13g2_buf_8 fanout2395 (.A(net2397),
    .X(net2395));
 sg13g2_buf_8 fanout2396 (.A(net2397),
    .X(net2396));
 sg13g2_buf_8 fanout2397 (.A(net2398),
    .X(net2397));
 sg13g2_buf_8 fanout2398 (.A(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2398));
 sg13g2_buf_8 fanout2399 (.A(net2400),
    .X(net2399));
 sg13g2_buf_8 fanout2400 (.A(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_nand2_1_A_Y ),
    .X(net2400));
 sg13g2_buf_8 fanout2401 (.A(net2406),
    .X(net2401));
 sg13g2_buf_8 fanout2402 (.A(net2406),
    .X(net2402));
 sg13g2_buf_8 fanout2403 (.A(net2406),
    .X(net2403));
 sg13g2_buf_1 fanout2404 (.A(net2405),
    .X(net2404));
 sg13g2_buf_8 fanout2405 (.A(net2406),
    .X(net2405));
 sg13g2_buf_8 fanout2406 (.A(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2406));
 sg13g2_buf_8 fanout2407 (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .X(net2407));
 sg13g2_buf_8 fanout2408 (.A(\i_snitch.pc_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .X(net2408));
 sg13g2_buf_8 fanout2409 (.A(net2410),
    .X(net2409));
 sg13g2_buf_8 fanout2410 (.A(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y ),
    .X(net2410));
 sg13g2_buf_8 fanout2411 (.A(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y ),
    .X(net2411));
 sg13g2_buf_8 fanout2412 (.A(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor3_1_A_C_sg13g2_nor2_1_B_Y ),
    .X(net2412));
 sg13g2_buf_8 fanout2413 (.A(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .X(net2413));
 sg13g2_buf_8 fanout2414 (.A(\i_snitch.i_snitch_regfile.mem[96]_sg13g2_dfrbpq_1_Q_D_sg13g2_o21ai_1_Y_A2 ),
    .X(net2414));
 sg13g2_buf_2 fanout2415 (.A(net2416),
    .X(net2415));
 sg13g2_buf_1 fanout2416 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2416));
 sg13g2_buf_2 fanout2417 (.A(net2418),
    .X(net2417));
 sg13g2_buf_1 fanout2418 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2418));
 sg13g2_buf_2 fanout2419 (.A(net2420),
    .X(net2419));
 sg13g2_buf_2 fanout2420 (.A(net2421),
    .X(net2420));
 sg13g2_buf_1 fanout2421 (.A(net2422),
    .X(net2421));
 sg13g2_buf_8 fanout2422 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2422));
 sg13g2_buf_8 fanout2423 (.A(net2428),
    .X(net2423));
 sg13g2_buf_8 fanout2424 (.A(net2428),
    .X(net2424));
 sg13g2_buf_8 fanout2425 (.A(net2427),
    .X(net2425));
 sg13g2_buf_8 fanout2426 (.A(net2427),
    .X(net2426));
 sg13g2_buf_8 fanout2427 (.A(net2428),
    .X(net2427));
 sg13g2_buf_8 fanout2428 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_or2_1_A_X ),
    .X(net2428));
 sg13g2_buf_8 fanout2429 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_and2_1_B_X_sg13g2_nor2_1_A_Y ),
    .X(net2429));
 sg13g2_buf_8 fanout2430 (.A(net2432),
    .X(net2430));
 sg13g2_buf_8 fanout2431 (.A(net2432),
    .X(net2431));
 sg13g2_buf_8 fanout2432 (.A(\i_snitch.sb_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2432));
 sg13g2_buf_8 fanout2433 (.A(net2435),
    .X(net2433));
 sg13g2_buf_8 fanout2434 (.A(net2435),
    .X(net2434));
 sg13g2_buf_8 fanout2435 (.A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2435));
 sg13g2_buf_8 fanout2436 (.A(net2438),
    .X(net2436));
 sg13g2_buf_8 fanout2437 (.A(net2438),
    .X(net2437));
 sg13g2_buf_8 fanout2438 (.A(\i_snitch.sb_d[7]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2438));
 sg13g2_buf_8 fanout2439 (.A(net2441),
    .X(net2439));
 sg13g2_buf_8 fanout2440 (.A(net2441),
    .X(net2440));
 sg13g2_buf_8 fanout2441 (.A(\i_snitch.sb_d[6]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2441));
 sg13g2_buf_8 fanout2442 (.A(net2444),
    .X(net2442));
 sg13g2_buf_8 fanout2443 (.A(net2444),
    .X(net2443));
 sg13g2_buf_8 fanout2444 (.A(\i_snitch.sb_d[5]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2444));
 sg13g2_buf_8 fanout2445 (.A(net2447),
    .X(net2445));
 sg13g2_buf_8 fanout2446 (.A(net2447),
    .X(net2446));
 sg13g2_buf_8 fanout2447 (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2447));
 sg13g2_buf_8 fanout2448 (.A(net2449),
    .X(net2448));
 sg13g2_buf_8 fanout2449 (.A(net2450),
    .X(net2449));
 sg13g2_buf_8 fanout2450 (.A(\i_snitch.sb_d[3]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_A_Y ),
    .X(net2450));
 sg13g2_buf_8 fanout2451 (.A(net2452),
    .X(net2451));
 sg13g2_buf_8 fanout2452 (.A(net2453),
    .X(net2452));
 sg13g2_buf_8 fanout2453 (.A(\i_snitch.sb_d[2]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2453));
 sg13g2_buf_8 fanout2454 (.A(net2455),
    .X(net2454));
 sg13g2_buf_8 fanout2455 (.A(net2456),
    .X(net2455));
 sg13g2_buf_8 fanout2456 (.A(\i_snitch.sb_d[1]_sg13g2_o21ai_1_Y_A1_sg13g2_nor3_1_B_Y ),
    .X(net2456));
 sg13g2_buf_8 fanout2457 (.A(net2459),
    .X(net2457));
 sg13g2_buf_8 fanout2458 (.A(net2459),
    .X(net2458));
 sg13g2_buf_8 fanout2459 (.A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2459));
 sg13g2_buf_8 fanout2460 (.A(net2462),
    .X(net2460));
 sg13g2_buf_8 fanout2461 (.A(net2462),
    .X(net2461));
 sg13g2_buf_8 fanout2462 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2462));
 sg13g2_buf_8 fanout2463 (.A(net2465),
    .X(net2463));
 sg13g2_buf_8 fanout2464 (.A(net2465),
    .X(net2464));
 sg13g2_buf_8 fanout2465 (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2465));
 sg13g2_buf_8 fanout2466 (.A(net2468),
    .X(net2466));
 sg13g2_buf_8 fanout2467 (.A(net2468),
    .X(net2467));
 sg13g2_buf_8 fanout2468 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2468));
 sg13g2_buf_8 fanout2469 (.A(net2471),
    .X(net2469));
 sg13g2_buf_8 fanout2470 (.A(net2471),
    .X(net2470));
 sg13g2_buf_8 fanout2471 (.A(\i_snitch.sb_d[11]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2471));
 sg13g2_buf_8 fanout2472 (.A(net2474),
    .X(net2472));
 sg13g2_buf_8 fanout2473 (.A(net2474),
    .X(net2473));
 sg13g2_buf_8 fanout2474 (.A(\i_snitch.sb_d[10]_sg13g2_o21ai_1_Y_A2_sg13g2_nor3_1_B_Y ),
    .X(net2474));
 sg13g2_buf_8 fanout2475 (.A(net2476),
    .X(net2475));
 sg13g2_buf_8 fanout2476 (.A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_a22oi_1_A2_Y ),
    .X(net2476));
 sg13g2_buf_8 fanout2477 (.A(net2478),
    .X(net2477));
 sg13g2_buf_8 fanout2478 (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .X(net2478));
 sg13g2_buf_8 fanout2479 (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y ),
    .X(net2479));
 sg13g2_buf_2 fanout2480 (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y ),
    .X(net2480));
 sg13g2_buf_8 fanout2481 (.A(net2483),
    .X(net2481));
 sg13g2_buf_1 fanout2482 (.A(net2483),
    .X(net2482));
 sg13g2_buf_2 fanout2483 (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B2_sg13g2_a221oi_1_A2_Y_sg13g2_nor2_1_A_Y ),
    .X(net2483));
 sg13g2_buf_8 fanout2484 (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .X(net2484));
 sg13g2_buf_8 fanout2485 (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_inv_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .X(net2485));
 sg13g2_buf_8 fanout2486 (.A(net2488),
    .X(net2486));
 sg13g2_buf_1 fanout2487 (.A(net2488),
    .X(net2487));
 sg13g2_buf_8 fanout2488 (.A(\i_snitch.i_snitch_lsu.handshake_pending_q_sg13g2_nor2_1_A_Y ),
    .X(net2488));
 sg13g2_buf_8 fanout2489 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ),
    .X(net2489));
 sg13g2_buf_8 fanout2490 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A_sg13g2_a22oi_1_Y_B2_sg13g2_o21ai_1_Y_A2_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ),
    .X(net2490));
 sg13g2_buf_8 fanout2491 (.A(net2492),
    .X(net2491));
 sg13g2_buf_8 fanout2492 (.A(net2493),
    .X(net2492));
 sg13g2_buf_8 fanout2493 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_o21ai_1_A2_Y ),
    .X(net2493));
 sg13g2_buf_8 fanout2494 (.A(net2497),
    .X(net2494));
 sg13g2_buf_8 fanout2495 (.A(net2497),
    .X(net2495));
 sg13g2_buf_8 fanout2496 (.A(net2497),
    .X(net2496));
 sg13g2_buf_8 fanout2497 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_o21ai_1_A2_Y ),
    .X(net2497));
 sg13g2_buf_8 fanout2498 (.A(net2502),
    .X(net2498));
 sg13g2_buf_8 fanout2499 (.A(net2502),
    .X(net2499));
 sg13g2_buf_8 fanout2500 (.A(net2501),
    .X(net2500));
 sg13g2_buf_8 fanout2501 (.A(net2502),
    .X(net2501));
 sg13g2_buf_8 fanout2502 (.A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_A1_sg13g2_nand2_1_A_Y ),
    .X(net2502));
 sg13g2_buf_8 fanout2503 (.A(net2505),
    .X(net2503));
 sg13g2_buf_1 fanout2504 (.A(net2505),
    .X(net2504));
 sg13g2_buf_8 fanout2505 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y ),
    .X(net2505));
 sg13g2_buf_8 fanout2506 (.A(net2507),
    .X(net2506));
 sg13g2_buf_8 fanout2507 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_or3_1_A_X_sg13g2_a22oi_1_B2_Y_sg13g2_nand3_1_C_Y ),
    .X(net2507));
 sg13g2_buf_8 fanout2508 (.A(net2511),
    .X(net2508));
 sg13g2_buf_2 fanout2509 (.A(net2511),
    .X(net2509));
 sg13g2_buf_8 fanout2510 (.A(net2511),
    .X(net2510));
 sg13g2_buf_8 fanout2511 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_nand2_1_B_Y ),
    .X(net2511));
 sg13g2_buf_8 fanout2512 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_and2_1_A_X_sg13g2_or4_1_C_X_sg13g2_and2_1_B_X ),
    .X(net2512));
 sg13g2_buf_8 fanout2513 (.A(net2514),
    .X(net2513));
 sg13g2_buf_8 fanout2514 (.A(\i_snitch.pc_d[1]_sg13g2_o21ai_1_Y_A2_sg13g2_a21oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_o21ai_1_A2_Y ),
    .X(net2514));
 sg13g2_buf_8 fanout2515 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y ),
    .X(net2515));
 sg13g2_buf_1 fanout2516 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_nor2_1_B_Y ),
    .X(net2516));
 sg13g2_buf_8 fanout2517 (.A(net2518),
    .X(net2517));
 sg13g2_buf_8 fanout2518 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X ),
    .X(net2518));
 sg13g2_buf_8 fanout2519 (.A(net2520),
    .X(net2519));
 sg13g2_buf_8 fanout2520 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y_sg13g2_and2_1_A_X ),
    .X(net2520));
 sg13g2_buf_8 fanout2521 (.A(\i_snitch.consec_pc[0]_sg13g2_a22oi_1_A1_Y ),
    .X(net2521));
 sg13g2_buf_8 fanout2522 (.A(\i_snitch.consec_pc[0]_sg13g2_a22oi_1_A1_Y ),
    .X(net2522));
 sg13g2_buf_8 fanout2523 (.A(net2529),
    .X(net2523));
 sg13g2_buf_2 fanout2524 (.A(net2529),
    .X(net2524));
 sg13g2_buf_8 fanout2525 (.A(net2529),
    .X(net2525));
 sg13g2_buf_1 fanout2526 (.A(net2529),
    .X(net2526));
 sg13g2_buf_8 fanout2527 (.A(net2528),
    .X(net2527));
 sg13g2_buf_8 fanout2528 (.A(net2529),
    .X(net2528));
 sg13g2_buf_8 fanout2529 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X_sg13g2_and2_1_A_X ),
    .X(net2529));
 sg13g2_buf_8 fanout2530 (.A(net2534),
    .X(net2530));
 sg13g2_buf_1 fanout2531 (.A(net2534),
    .X(net2531));
 sg13g2_buf_8 fanout2532 (.A(net2534),
    .X(net2532));
 sg13g2_buf_8 fanout2533 (.A(net2534),
    .X(net2533));
 sg13g2_buf_8 fanout2534 (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_nand4_1_D_B_sg13g2_nand2_1_B_Y_sg13g2_nand2_1_B_Y ),
    .X(net2534));
 sg13g2_buf_16 fanout2535 (.X(net2535),
    .A(net2536));
 sg13g2_buf_16 fanout2536 (.X(net2536),
    .A(net2537));
 sg13g2_buf_16 fanout2537 (.X(net2537),
    .A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nand2b_1_B_A_N_sg13g2_nor3_1_C_B_sg13g2_and3_1_A_X ));
 sg13g2_buf_8 fanout2538 (.A(net2539),
    .X(net2538));
 sg13g2_buf_8 fanout2539 (.A(\i_snitch.pc_d[9]_sg13g2_o21ai_1_Y_A2_sg13g2_a22oi_1_Y_A2_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_o21ai_1_Y_A2_sg13g2_mux2_1_X_A1_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A_sg13g2_nor2_1_B_Y ),
    .X(net2539));
 sg13g2_buf_8 fanout2540 (.A(net2541),
    .X(net2540));
 sg13g2_buf_8 fanout2541 (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_nand2_1_A_Y ),
    .X(net2541));
 sg13g2_buf_8 fanout2542 (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X ),
    .X(net2542));
 sg13g2_buf_8 fanout2543 (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_A1_sg13g2_and2_1_X_A_sg13g2_and2_1_A_X ),
    .X(net2543));
 sg13g2_buf_8 fanout2544 (.A(net2545),
    .X(net2544));
 sg13g2_buf_8 fanout2545 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y ),
    .X(net2545));
 sg13g2_buf_8 fanout2546 (.A(net2547),
    .X(net2546));
 sg13g2_buf_8 fanout2547 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_B_sg13g2_nor4_1_Y_B_sg13g2_or2_1_B_X_sg13g2_nand2b_1_A_N_Y ),
    .X(net2547));
 sg13g2_buf_8 fanout2548 (.A(\i_snitch.i_snitch_regfile.mem[438]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(net2548));
 sg13g2_buf_8 fanout2549 (.A(net2550),
    .X(net2549));
 sg13g2_buf_8 fanout2550 (.A(net2553),
    .X(net2550));
 sg13g2_buf_8 fanout2551 (.A(net2552),
    .X(net2551));
 sg13g2_buf_8 fanout2552 (.A(net2553),
    .X(net2552));
 sg13g2_buf_8 fanout2553 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_Y_sg13g2_and4_1_D_X_sg13g2_nand3_1_C_A_sg13g2_nand3b_1_C_Y ),
    .X(net2553));
 sg13g2_buf_8 fanout2554 (.A(net2556),
    .X(net2554));
 sg13g2_buf_1 fanout2555 (.A(net2556),
    .X(net2555));
 sg13g2_buf_8 fanout2556 (.A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net2556));
 sg13g2_buf_8 fanout2557 (.A(net2559),
    .X(net2557));
 sg13g2_buf_1 fanout2558 (.A(net2559),
    .X(net2558));
 sg13g2_buf_1 fanout2559 (.A(net2560),
    .X(net2559));
 sg13g2_buf_8 fanout2560 (.A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net2560));
 sg13g2_buf_8 fanout2561 (.A(net2563),
    .X(net2561));
 sg13g2_buf_1 fanout2562 (.A(net88),
    .X(net2562));
 sg13g2_buf_8 fanout2563 (.A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ),
    .X(net2563));
 sg13g2_buf_8 fanout2564 (.A(net2568),
    .X(net2564));
 sg13g2_buf_8 fanout2565 (.A(net2567),
    .X(net2565));
 sg13g2_buf_8 fanout2566 (.A(net2567),
    .X(net2566));
 sg13g2_buf_8 fanout2567 (.A(net2568),
    .X(net2567));
 sg13g2_buf_8 fanout2568 (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21oi_1_B1_Y ),
    .X(net2568));
 sg13g2_buf_8 fanout2569 (.A(net2570),
    .X(net2569));
 sg13g2_buf_8 fanout2570 (.A(\i_snitch.i_snitch_regfile.mem[63]_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_a221oi_1_B2_Y_sg13g2_mux2_1_S_A0_sg13g2_a21o_1_B1_X ),
    .X(net2570));
 sg13g2_buf_8 fanout2571 (.A(net2575),
    .X(net2571));
 sg13g2_buf_8 fanout2572 (.A(net2574),
    .X(net2572));
 sg13g2_buf_1 fanout2573 (.A(net2574),
    .X(net2573));
 sg13g2_buf_8 fanout2574 (.A(net2575),
    .X(net2574));
 sg13g2_buf_2 fanout2575 (.A(net2576),
    .X(net2575));
 sg13g2_buf_8 fanout2576 (.A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net2576));
 sg13g2_buf_8 fanout2577 (.A(net2578),
    .X(net2577));
 sg13g2_buf_8 fanout2578 (.A(net2579),
    .X(net2578));
 sg13g2_buf_8 fanout2579 (.A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand2b_1_A_N_Y ),
    .X(net2579));
 sg13g2_buf_2 fanout2580 (.A(net2583),
    .X(net2580));
 sg13g2_buf_8 fanout2581 (.A(net2583),
    .X(net2581));
 sg13g2_buf_1 fanout2582 (.A(net2583),
    .X(net2582));
 sg13g2_buf_8 fanout2583 (.A(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2583));
 sg13g2_buf_8 fanout2584 (.A(net2585),
    .X(net2584));
 sg13g2_buf_2 fanout2585 (.A(net2588),
    .X(net2585));
 sg13g2_buf_8 fanout2586 (.A(net2587),
    .X(net2586));
 sg13g2_buf_8 fanout2587 (.A(net2588),
    .X(net2587));
 sg13g2_buf_1 fanout2588 (.A(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2588));
 sg13g2_buf_8 fanout2589 (.A(\i_snitch.i_snitch_regfile.mem[35]_sg13g2_a22oi_1_A1_Y_sg13g2_a221oi_1_B1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2589));
 sg13g2_buf_8 fanout2590 (.A(net2591),
    .X(net2590));
 sg13g2_buf_2 fanout2591 (.A(net2592),
    .X(net2591));
 sg13g2_buf_8 fanout2592 (.A(net2593),
    .X(net2592));
 sg13g2_buf_8 fanout2593 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand3_1_C_Y ),
    .X(net2593));
 sg13g2_buf_8 fanout2594 (.A(net2595),
    .X(net2594));
 sg13g2_buf_1 fanout2595 (.A(net2598),
    .X(net2595));
 sg13g2_buf_2 fanout2596 (.A(net2597),
    .X(net2596));
 sg13g2_buf_1 fanout2597 (.A(net2598),
    .X(net2597));
 sg13g2_buf_1 fanout2598 (.A(net2599),
    .X(net2598));
 sg13g2_buf_8 fanout2599 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_Y_sg13g2_and3_1_C_X ),
    .X(net2599));
 sg13g2_buf_8 fanout2600 (.A(net2602),
    .X(net2600));
 sg13g2_buf_1 fanout2601 (.A(net2602),
    .X(net2601));
 sg13g2_buf_8 fanout2602 (.A(net2603),
    .X(net2602));
 sg13g2_buf_8 fanout2603 (.A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net2603));
 sg13g2_buf_2 fanout2604 (.A(net2605),
    .X(net2604));
 sg13g2_buf_1 fanout2605 (.A(net2606),
    .X(net2605));
 sg13g2_buf_1 fanout2606 (.A(net2607),
    .X(net2606));
 sg13g2_buf_1 fanout2607 (.A(net65),
    .X(net2607));
 sg13g2_buf_16 fanout2608 (.X(net2608),
    .A(net2609));
 sg13g2_buf_8 fanout2609 (.A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nand2b_1_A_N_Y ),
    .X(net2609));
 sg13g2_buf_8 fanout2610 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_or4_1_C_X ),
    .X(net2610));
 sg13g2_buf_8 fanout2611 (.A(net2612),
    .X(net2611));
 sg13g2_buf_8 fanout2612 (.A(net2615),
    .X(net2612));
 sg13g2_buf_8 fanout2613 (.A(net2615),
    .X(net2613));
 sg13g2_buf_1 fanout2614 (.A(net2615),
    .X(net2614));
 sg13g2_buf_8 fanout2615 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_Y_sg13g2_a21o_1_A2_X_sg13g2_or4_1_B_X_sg13g2_nor4_1_C_Y ),
    .X(net2615));
 sg13g2_buf_8 fanout2616 (.A(net2618),
    .X(net2616));
 sg13g2_buf_8 fanout2617 (.A(net2618),
    .X(net2617));
 sg13g2_buf_8 fanout2618 (.A(net2620),
    .X(net2618));
 sg13g2_buf_8 fanout2619 (.A(net2620),
    .X(net2619));
 sg13g2_buf_8 fanout2620 (.A(net2625),
    .X(net2620));
 sg13g2_buf_8 fanout2621 (.A(net2625),
    .X(net2621));
 sg13g2_buf_8 fanout2622 (.A(net2625),
    .X(net2622));
 sg13g2_buf_8 fanout2623 (.A(net2624),
    .X(net2623));
 sg13g2_buf_8 fanout2624 (.A(net2625),
    .X(net2624));
 sg13g2_buf_8 fanout2625 (.A(target_sel_q_sg13g2_nor2_1_A_B_sg13g2_nor2_1_Y_B_sg13g2_nand3b_1_B_Y),
    .X(net2625));
 sg13g2_buf_8 fanout2626 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_or2_1_B_X ),
    .X(net2626));
 sg13g2_buf_8 fanout2627 (.A(net2628),
    .X(net2627));
 sg13g2_buf_8 fanout2628 (.A(net2630),
    .X(net2628));
 sg13g2_buf_8 fanout2629 (.A(net2630),
    .X(net2629));
 sg13g2_buf_8 fanout2630 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_or2_1_A_X_sg13g2_a221oi_1_A2_B1_sg13g2_nor2_1_B_Y ),
    .X(net2630));
 sg13g2_buf_8 fanout2631 (.A(net2632),
    .X(net2631));
 sg13g2_buf_8 fanout2632 (.A(net2633),
    .X(net2632));
 sg13g2_buf_8 fanout2633 (.A(\i_snitch.i_snitch_regfile.mem[40]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a221oi_1_B2_C1_sg13g2_and2_1_X_B_sg13g2_nand2_1_B_Y ),
    .X(net2633));
 sg13g2_buf_8 fanout2634 (.A(net2636),
    .X(net2634));
 sg13g2_buf_8 fanout2635 (.A(net2636),
    .X(net2635));
 sg13g2_buf_8 fanout2636 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ),
    .X(net2636));
 sg13g2_buf_8 fanout2637 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X_sg13g2_nand2_1_A_Y ),
    .X(net2637));
 sg13g2_buf_8 fanout2638 (.A(net2640),
    .X(net2638));
 sg13g2_buf_8 fanout2639 (.A(net2640),
    .X(net2639));
 sg13g2_buf_8 fanout2640 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .X(net2640));
 sg13g2_buf_8 fanout2641 (.A(net2642),
    .X(net2641));
 sg13g2_buf_8 fanout2642 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_Y_sg13g2_nor3_1_C_Y ),
    .X(net2642));
 sg13g2_buf_8 fanout2643 (.A(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .X(net2643));
 sg13g2_buf_8 fanout2644 (.A(\data_pdata[8]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .X(net2644));
 sg13g2_buf_8 fanout2645 (.A(net2646),
    .X(net2645));
 sg13g2_buf_8 fanout2646 (.A(\data_pdata[31]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2646));
 sg13g2_buf_8 fanout2647 (.A(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2647));
 sg13g2_buf_2 fanout2648 (.A(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2648));
 sg13g2_buf_8 fanout2649 (.A(net2650),
    .X(net2649));
 sg13g2_buf_8 fanout2650 (.A(\data_pdata[30]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2650));
 sg13g2_buf_8 fanout2651 (.A(net2652),
    .X(net2651));
 sg13g2_buf_8 fanout2652 (.A(\data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2652));
 sg13g2_buf_8 fanout2653 (.A(net2654),
    .X(net2653));
 sg13g2_buf_8 fanout2654 (.A(\data_pdata[29]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2654));
 sg13g2_buf_8 fanout2655 (.A(net2656),
    .X(net2655));
 sg13g2_buf_8 fanout2656 (.A(\data_pdata[28]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2656));
 sg13g2_buf_8 fanout2657 (.A(net2658),
    .X(net2657));
 sg13g2_buf_8 fanout2658 (.A(\data_pdata[27]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2658));
 sg13g2_buf_8 fanout2659 (.A(net2660),
    .X(net2659));
 sg13g2_buf_8 fanout2660 (.A(\data_pdata[26]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2660));
 sg13g2_buf_8 fanout2661 (.A(net2662),
    .X(net2661));
 sg13g2_buf_8 fanout2662 (.A(\data_pdata[25]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2662));
 sg13g2_buf_8 fanout2663 (.A(\data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2663));
 sg13g2_buf_8 fanout2664 (.A(\data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2664));
 sg13g2_buf_8 fanout2665 (.A(net2666),
    .X(net2665));
 sg13g2_buf_8 fanout2666 (.A(\data_pdata[24]_sg13g2_nand2b_1_B_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2666));
 sg13g2_buf_8 fanout2667 (.A(net2668),
    .X(net2667));
 sg13g2_buf_8 fanout2668 (.A(\data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2668));
 sg13g2_buf_8 fanout2669 (.A(net2670),
    .X(net2669));
 sg13g2_buf_8 fanout2670 (.A(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_inv_1_A_Y_sg13g2_o21ai_1_A1_Y ),
    .X(net2670));
 sg13g2_buf_8 fanout2671 (.A(net2672),
    .X(net2671));
 sg13g2_buf_8 fanout2672 (.A(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .X(net2672));
 sg13g2_buf_8 fanout2673 (.A(net2674),
    .X(net2673));
 sg13g2_buf_8 fanout2674 (.A(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .X(net2674));
 sg13g2_buf_8 fanout2675 (.A(net2676),
    .X(net2675));
 sg13g2_buf_8 fanout2676 (.A(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_nand3b_1_C_Y_sg13g2_nand2_1_B_Y ),
    .X(net2676));
 sg13g2_buf_8 fanout2677 (.A(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .X(net2677));
 sg13g2_buf_8 fanout2678 (.A(\data_pdata[15]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_B1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .X(net2678));
 sg13g2_buf_8 fanout2679 (.A(net2680),
    .X(net2679));
 sg13g2_buf_8 fanout2680 (.A(\data_pdata[11]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21oi_1_A2_Y_sg13g2_inv_1_A_Y ),
    .X(net2680));
 sg13g2_buf_8 fanout2681 (.A(net2682),
    .X(net2681));
 sg13g2_buf_2 fanout2682 (.A(net2683),
    .X(net2682));
 sg13g2_buf_2 fanout2683 (.A(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_nand4_1_A_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net2683));
 sg13g2_buf_8 fanout2684 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_nor2_1_A_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2684));
 sg13g2_buf_8 fanout2685 (.A(net2686),
    .X(net2685));
 sg13g2_buf_8 fanout2686 (.A(\data_pdata[9]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2686));
 sg13g2_buf_8 fanout2687 (.A(\data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2687));
 sg13g2_buf_8 fanout2688 (.A(\data_pdata[14]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2688));
 sg13g2_buf_8 fanout2689 (.A(\data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2689));
 sg13g2_buf_8 fanout2690 (.A(\data_pdata[13]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2690));
 sg13g2_buf_8 fanout2691 (.A(net2692),
    .X(net2691));
 sg13g2_buf_8 fanout2692 (.A(\data_pdata[12]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2692));
 sg13g2_buf_8 fanout2693 (.A(net2694),
    .X(net2693));
 sg13g2_buf_8 fanout2694 (.A(\data_pdata[10]_sg13g2_nand2b_1_B_Y_sg13g2_a22oi_1_A1_Y_sg13g2_a21o_1_A2_X ),
    .X(net2694));
 sg13g2_buf_8 fanout2695 (.A(net2698),
    .X(net2695));
 sg13g2_buf_8 fanout2696 (.A(net2698),
    .X(net2696));
 sg13g2_buf_2 fanout2697 (.A(net2698),
    .X(net2697));
 sg13g2_buf_8 fanout2698 (.A(\i_snitch.pc_d[6]_sg13g2_mux2_1_X_A1_sg13g2_a21o_1_X_A2_sg13g2_xor2_1_X_A_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_B_sg13g2_nand4_1_A_C_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_a21o_1_B1_X ),
    .X(net2698));
 sg13g2_buf_8 fanout2699 (.A(net2703),
    .X(net2699));
 sg13g2_buf_8 fanout2700 (.A(net2702),
    .X(net2700));
 sg13g2_buf_1 fanout2701 (.A(net2702),
    .X(net2701));
 sg13g2_buf_2 fanout2702 (.A(net2703),
    .X(net2702));
 sg13g2_buf_8 fanout2703 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X ),
    .X(net2703));
 sg13g2_buf_8 fanout2704 (.A(net2705),
    .X(net2704));
 sg13g2_buf_8 fanout2705 (.A(net2708),
    .X(net2705));
 sg13g2_buf_8 fanout2706 (.A(net2707),
    .X(net2706));
 sg13g2_buf_8 fanout2707 (.A(net2708),
    .X(net2707));
 sg13g2_buf_8 fanout2708 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_X ),
    .X(net2708));
 sg13g2_buf_8 fanout2709 (.A(net2710),
    .X(net2709));
 sg13g2_buf_1 fanout2710 (.A(net2711),
    .X(net2710));
 sg13g2_buf_2 fanout2711 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X ),
    .X(net2711));
 sg13g2_buf_8 fanout2712 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X ),
    .X(net2712));
 sg13g2_buf_1 fanout2713 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_X ),
    .X(net2713));
 sg13g2_buf_8 fanout2714 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_nand2_1_A_Y_sg13g2_nor2_1_B_Y ),
    .X(net2714));
 sg13g2_buf_8 fanout2715 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net2715));
 sg13g2_buf_8 fanout2716 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand2b_1_A_N_Y ),
    .X(net2716));
 sg13g2_buf_8 fanout2717 (.A(net2718),
    .X(net2717));
 sg13g2_buf_8 fanout2718 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net2718));
 sg13g2_buf_8 fanout2719 (.A(net2721),
    .X(net2719));
 sg13g2_buf_8 fanout2720 (.A(net2721),
    .X(net2720));
 sg13g2_buf_8 fanout2721 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X ),
    .X(net2721));
 sg13g2_buf_8 fanout2722 (.A(net2726),
    .X(net2722));
 sg13g2_buf_1 fanout2723 (.A(net2726),
    .X(net2723));
 sg13g2_buf_8 fanout2724 (.A(net2726),
    .X(net2724));
 sg13g2_buf_8 fanout2725 (.A(net2726),
    .X(net2725));
 sg13g2_buf_8 fanout2726 (.A(net97),
    .X(net2726));
 sg13g2_buf_8 fanout2727 (.A(net2729),
    .X(net2727));
 sg13g2_buf_8 fanout2728 (.A(net2729),
    .X(net2728));
 sg13g2_buf_8 fanout2729 (.A(net2730),
    .X(net2729));
 sg13g2_buf_8 fanout2730 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y ),
    .X(net2730));
 sg13g2_buf_8 fanout2731 (.A(net2732),
    .X(net2731));
 sg13g2_buf_8 fanout2732 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y ),
    .X(net2732));
 sg13g2_buf_8 fanout2733 (.A(net2734),
    .X(net2733));
 sg13g2_buf_8 fanout2734 (.A(net2737),
    .X(net2734));
 sg13g2_buf_2 fanout2735 (.A(net2736),
    .X(net2735));
 sg13g2_buf_1 fanout2736 (.A(net2737),
    .X(net2736));
 sg13g2_buf_8 fanout2737 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_nor2_1_B_A_sg13g2_nand2b_1_B_Y ),
    .X(net2737));
 sg13g2_buf_8 fanout2738 (.A(net2740),
    .X(net2738));
 sg13g2_buf_8 fanout2739 (.A(net2740),
    .X(net2739));
 sg13g2_buf_8 fanout2740 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2740));
 sg13g2_buf_8 fanout2741 (.A(net2743),
    .X(net2741));
 sg13g2_buf_8 fanout2742 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2742));
 sg13g2_buf_8 fanout2743 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1_sg13g2_o21ai_1_Y_A1_sg13g2_nor2_1_A_Y ),
    .X(net2743));
 sg13g2_buf_8 fanout2744 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ),
    .X(net2744));
 sg13g2_buf_8 fanout2745 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y ),
    .X(net2745));
 sg13g2_buf_1 fanout2746 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y ),
    .X(net2746));
 sg13g2_buf_8 fanout2747 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21oi_1_B1_Y ),
    .X(net2747));
 sg13g2_buf_8 fanout2748 (.A(net2749),
    .X(net2748));
 sg13g2_buf_8 fanout2749 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_D_sg13g2_or4_1_X_C_sg13g2_a21o_1_B1_X ),
    .X(net2749));
 sg13g2_buf_8 fanout2750 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand4_1_B_A_sg13g2_nor3_1_B_A_sg13g2_nor3_1_A_Y_sg13g2_a22oi_1_A2_Y ),
    .X(net2750));
 sg13g2_buf_8 fanout2751 (.A(net2754),
    .X(net2751));
 sg13g2_buf_2 fanout2752 (.A(net2754),
    .X(net2752));
 sg13g2_buf_8 fanout2753 (.A(net2754),
    .X(net2753));
 sg13g2_buf_8 fanout2754 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nor2_1_B_Y ),
    .X(net2754));
 sg13g2_buf_8 fanout2755 (.A(net2756),
    .X(net2755));
 sg13g2_buf_2 fanout2756 (.A(net2763),
    .X(net2756));
 sg13g2_buf_8 fanout2757 (.A(net2758),
    .X(net2757));
 sg13g2_buf_8 fanout2758 (.A(net2763),
    .X(net2758));
 sg13g2_buf_8 fanout2759 (.A(net2760),
    .X(net2759));
 sg13g2_buf_8 fanout2760 (.A(net2763),
    .X(net2760));
 sg13g2_buf_8 fanout2761 (.A(net2763),
    .X(net2761));
 sg13g2_buf_2 fanout2762 (.A(net2763),
    .X(net2762));
 sg13g2_buf_8 fanout2763 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_nand4_1_D_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2763));
 sg13g2_buf_8 fanout2764 (.A(net2766),
    .X(net2764));
 sg13g2_buf_1 fanout2765 (.A(net2766),
    .X(net2765));
 sg13g2_buf_1 fanout2766 (.A(net2770),
    .X(net2766));
 sg13g2_buf_8 fanout2767 (.A(net2770),
    .X(net2767));
 sg13g2_buf_8 fanout2768 (.A(net2770),
    .X(net2768));
 sg13g2_buf_8 fanout2769 (.A(net2770),
    .X(net2769));
 sg13g2_buf_8 fanout2770 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_2_X),
    .X(net2770));
 sg13g2_buf_8 fanout2771 (.A(net2772),
    .X(net2771));
 sg13g2_buf_8 fanout2772 (.A(net2773),
    .X(net2772));
 sg13g2_buf_8 fanout2773 (.A(net2776),
    .X(net2773));
 sg13g2_buf_8 fanout2774 (.A(net2776),
    .X(net2774));
 sg13g2_buf_8 fanout2775 (.A(net2776),
    .X(net2775));
 sg13g2_buf_8 fanout2776 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_1_X),
    .X(net2776));
 sg13g2_buf_8 fanout2777 (.A(net2778),
    .X(net2777));
 sg13g2_buf_8 fanout2778 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X),
    .X(net2778));
 sg13g2_buf_8 fanout2779 (.A(net2781),
    .X(net2779));
 sg13g2_buf_8 fanout2780 (.A(net2781),
    .X(net2780));
 sg13g2_buf_8 fanout2781 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_A_X),
    .X(net2781));
 sg13g2_buf_8 fanout2782 (.A(net2783),
    .X(net2782));
 sg13g2_buf_8 fanout2783 (.A(net2784),
    .X(net2783));
 sg13g2_buf_8 fanout2784 (.A(net2785),
    .X(net2784));
 sg13g2_buf_8 fanout2785 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X),
    .X(net2785));
 sg13g2_buf_8 fanout2786 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X),
    .X(net2786));
 sg13g2_buf_8 fanout2787 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_B_X),
    .X(net2787));
 sg13g2_buf_8 fanout2788 (.A(net2789),
    .X(net2788));
 sg13g2_buf_8 fanout2789 (.A(net2790),
    .X(net2789));
 sg13g2_buf_8 fanout2790 (.A(net2793),
    .X(net2790));
 sg13g2_buf_8 fanout2791 (.A(net2792),
    .X(net2791));
 sg13g2_buf_8 fanout2792 (.A(net2793),
    .X(net2792));
 sg13g2_buf_8 fanout2793 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_1_X),
    .X(net2793));
 sg13g2_buf_8 fanout2794 (.A(net2799),
    .X(net2794));
 sg13g2_buf_8 fanout2795 (.A(net2799),
    .X(net2795));
 sg13g2_buf_8 fanout2796 (.A(net2799),
    .X(net2796));
 sg13g2_buf_1 fanout2797 (.A(net2798),
    .X(net2797));
 sg13g2_buf_8 fanout2798 (.A(net2799),
    .X(net2798));
 sg13g2_buf_8 fanout2799 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y_sg13g2_and2_1_B_X_sg13g2_and2_1_A_X),
    .X(net2799));
 sg13g2_buf_8 fanout2800 (.A(net2801),
    .X(net2800));
 sg13g2_buf_8 fanout2801 (.A(net2802),
    .X(net2801));
 sg13g2_buf_8 fanout2802 (.A(net2809),
    .X(net2802));
 sg13g2_buf_2 fanout2803 (.A(net2809),
    .X(net2803));
 sg13g2_buf_8 fanout2804 (.A(net2809),
    .X(net2804));
 sg13g2_buf_1 fanout2805 (.A(net2809),
    .X(net2805));
 sg13g2_buf_8 fanout2806 (.A(net2807),
    .X(net2806));
 sg13g2_buf_8 fanout2807 (.A(net2808),
    .X(net2807));
 sg13g2_buf_8 fanout2808 (.A(net2809),
    .X(net2808));
 sg13g2_buf_8 fanout2809 (.A(\i_snitch.i_snitch_regfile.mem[98]_sg13g2_nor2_1_A_B ),
    .X(net2809));
 sg13g2_buf_8 fanout2810 (.A(net2813),
    .X(net2810));
 sg13g2_buf_8 fanout2811 (.A(net2813),
    .X(net2811));
 sg13g2_buf_8 fanout2812 (.A(net2813),
    .X(net2812));
 sg13g2_buf_8 fanout2813 (.A(\i_snitch.i_snitch_regfile.mem[420]_sg13g2_o21ai_1_A1_A2 ),
    .X(net2813));
 sg13g2_buf_8 fanout2814 (.A(\i_snitch.i_snitch_regfile.mem[259]_sg13g2_o21ai_1_A1_A2 ),
    .X(net2814));
 sg13g2_buf_8 fanout2815 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X_sg13g2_and4_1_D_X ),
    .X(net2815));
 sg13g2_buf_8 fanout2816 (.A(net2818),
    .X(net2816));
 sg13g2_buf_2 fanout2817 (.A(net2818),
    .X(net2817));
 sg13g2_buf_8 fanout2818 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y ),
    .X(net2818));
 sg13g2_buf_8 fanout2819 (.A(net2820),
    .X(net2819));
 sg13g2_buf_8 fanout2820 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y_sg13g2_nand2_1_A_1_Y ),
    .X(net2820));
 sg13g2_buf_8 fanout2821 (.A(net2823),
    .X(net2821));
 sg13g2_buf_8 fanout2822 (.A(net2823),
    .X(net2822));
 sg13g2_buf_8 fanout2823 (.A(\i_snitch.i_snitch_regfile.mem[53]_sg13g2_a21oi_1_A1_B1 ),
    .X(net2823));
 sg13g2_buf_8 fanout2824 (.A(net2825),
    .X(net2824));
 sg13g2_buf_8 fanout2825 (.A(net2826),
    .X(net2825));
 sg13g2_buf_8 fanout2826 (.A(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_A2 ),
    .X(net2826));
 sg13g2_buf_8 fanout2827 (.A(net2830),
    .X(net2827));
 sg13g2_buf_8 fanout2828 (.A(net2829),
    .X(net2828));
 sg13g2_buf_8 fanout2829 (.A(net2830),
    .X(net2829));
 sg13g2_buf_8 fanout2830 (.A(\i_snitch.i_snitch_regfile.mem[36]_sg13g2_a22oi_1_A1_A2 ),
    .X(net2830));
 sg13g2_buf_8 fanout2831 (.A(net2832),
    .X(net2831));
 sg13g2_buf_8 fanout2832 (.A(net2833),
    .X(net2832));
 sg13g2_buf_8 fanout2833 (.A(\i_snitch.i_snitch_regfile.mem[97]_sg13g2_o21ai_1_A1_B1 ),
    .X(net2833));
 sg13g2_buf_8 fanout2834 (.A(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_B1 ),
    .X(net2834));
 sg13g2_buf_8 fanout2835 (.A(\i_snitch.i_snitch_regfile.mem[94]_sg13g2_a21oi_1_A1_B1 ),
    .X(net2835));
 sg13g2_buf_8 fanout2836 (.A(net2837),
    .X(net2836));
 sg13g2_buf_8 fanout2837 (.A(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A ),
    .X(net2837));
 sg13g2_buf_8 fanout2838 (.A(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A ),
    .X(net2838));
 sg13g2_buf_8 fanout2839 (.A(\i_snitch.i_snitch_regfile.mem[128]_sg13g2_mux4_1_A0_1_X_sg13g2_nor2_1_B_A ),
    .X(net2839));
 sg13g2_buf_8 fanout2840 (.A(net2841),
    .X(net2840));
 sg13g2_buf_8 fanout2841 (.A(net2842),
    .X(net2841));
 sg13g2_buf_8 fanout2842 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y ),
    .X(net2842));
 sg13g2_buf_8 fanout2843 (.A(net2847),
    .X(net2843));
 sg13g2_buf_8 fanout2844 (.A(net2847),
    .X(net2844));
 sg13g2_buf_8 fanout2845 (.A(net2846),
    .X(net2845));
 sg13g2_buf_8 fanout2846 (.A(net2847),
    .X(net2846));
 sg13g2_buf_8 fanout2847 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y_sg13g2_nor2_1_B_Y ),
    .X(net2847));
 sg13g2_buf_8 fanout2848 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a22oi_1_A1_Y_sg13g2_nand2_1_B_Y ),
    .X(net2848));
 sg13g2_buf_8 fanout2849 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X ),
    .X(net2849));
 sg13g2_buf_1 fanout2850 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X ),
    .X(net2850));
 sg13g2_buf_8 fanout2851 (.A(net2853),
    .X(net2851));
 sg13g2_buf_2 fanout2852 (.A(net2853),
    .X(net2852));
 sg13g2_buf_8 fanout2853 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and2_1_B_X ),
    .X(net2853));
 sg13g2_buf_8 fanout2854 (.A(net2856),
    .X(net2854));
 sg13g2_buf_8 fanout2855 (.A(net2856),
    .X(net2855));
 sg13g2_buf_8 fanout2856 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y),
    .X(net2856));
 sg13g2_buf_8 fanout2857 (.A(net2859),
    .X(net2857));
 sg13g2_buf_8 fanout2858 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y),
    .X(net2858));
 sg13g2_buf_8 fanout2859 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand3_1_C_Y_sg13g2_nor2_1_A_Y),
    .X(net2859));
 sg13g2_buf_8 fanout2860 (.A(net2861),
    .X(net2860));
 sg13g2_buf_8 fanout2861 (.A(net2865),
    .X(net2861));
 sg13g2_buf_8 fanout2862 (.A(net2864),
    .X(net2862));
 sg13g2_buf_8 fanout2863 (.A(net2864),
    .X(net2863));
 sg13g2_buf_8 fanout2864 (.A(net2865),
    .X(net2864));
 sg13g2_buf_8 fanout2865 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_nand2_1_B_Y_sg13g2_nor3_1_B_Y),
    .X(net2865));
 sg13g2_buf_8 fanout2866 (.A(net2867),
    .X(net2866));
 sg13g2_buf_8 fanout2867 (.A(net2868),
    .X(net2867));
 sg13g2_buf_8 fanout2868 (.A(net2869),
    .X(net2868));
 sg13g2_buf_8 fanout2869 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X),
    .X(net2869));
 sg13g2_buf_8 fanout2870 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X),
    .X(net2870));
 sg13g2_buf_8 fanout2871 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_B_X),
    .X(net2871));
 sg13g2_buf_8 fanout2872 (.A(net2873),
    .X(net2872));
 sg13g2_buf_8 fanout2873 (.A(net2874),
    .X(net2873));
 sg13g2_buf_8 fanout2874 (.A(net2877),
    .X(net2874));
 sg13g2_buf_8 fanout2875 (.A(net2877),
    .X(net2875));
 sg13g2_buf_8 fanout2876 (.A(net2877),
    .X(net2876));
 sg13g2_buf_8 fanout2877 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_1_X),
    .X(net2877));
 sg13g2_buf_8 fanout2878 (.A(net2884),
    .X(net2878));
 sg13g2_buf_8 fanout2879 (.A(net2880),
    .X(net2879));
 sg13g2_buf_8 fanout2880 (.A(net2884),
    .X(net2880));
 sg13g2_buf_8 fanout2881 (.A(net2883),
    .X(net2881));
 sg13g2_buf_8 fanout2882 (.A(net2883),
    .X(net2882));
 sg13g2_buf_8 fanout2883 (.A(net2884),
    .X(net2883));
 sg13g2_buf_8 fanout2884 (.A(data_pvalid_sg13g2_nor2b_1_B_N_Y_sg13g2_and3_1_C_X_sg13g2_and2_1_A_X),
    .X(net2884));
 sg13g2_buf_8 fanout2885 (.A(net2886),
    .X(net2885));
 sg13g2_buf_8 fanout2886 (.A(net2887),
    .X(net2886));
 sg13g2_buf_8 fanout2887 (.A(net2890),
    .X(net2887));
 sg13g2_buf_8 fanout2888 (.A(net2889),
    .X(net2888));
 sg13g2_buf_8 fanout2889 (.A(net2890),
    .X(net2889));
 sg13g2_buf_8 fanout2890 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_1_X),
    .X(net2890));
 sg13g2_buf_8 fanout2891 (.A(net2896),
    .X(net2891));
 sg13g2_buf_8 fanout2892 (.A(net2896),
    .X(net2892));
 sg13g2_buf_8 fanout2893 (.A(net2894),
    .X(net2893));
 sg13g2_buf_8 fanout2894 (.A(net2896),
    .X(net2894));
 sg13g2_buf_8 fanout2895 (.A(net2896),
    .X(net2895));
 sg13g2_buf_8 fanout2896 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor3_1_C_Y_sg13g2_and2_1_A_X),
    .X(net2896));
 sg13g2_buf_8 fanout2897 (.A(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2897));
 sg13g2_buf_8 fanout2898 (.A(\data_pdata[31]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2898));
 sg13g2_buf_8 fanout2899 (.A(net2900),
    .X(net2899));
 sg13g2_buf_8 fanout2900 (.A(\data_pdata[30]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2900));
 sg13g2_buf_8 fanout2901 (.A(net2902),
    .X(net2901));
 sg13g2_buf_8 fanout2902 (.A(\data_pdata[25]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2902));
 sg13g2_buf_8 fanout2903 (.A(\data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2903));
 sg13g2_buf_8 fanout2904 (.A(\data_pdata[24]_sg13g2_a21oi_1_A2_Y_sg13g2_a21oi_1_A2_Y ),
    .X(net2904));
 sg13g2_buf_8 fanout2905 (.A(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2905));
 sg13g2_buf_8 fanout2906 (.A(\data_pdata[21]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2906));
 sg13g2_buf_8 fanout2907 (.A(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2907));
 sg13g2_buf_8 fanout2908 (.A(\data_pdata[20]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2908));
 sg13g2_buf_8 fanout2909 (.A(net2910),
    .X(net2909));
 sg13g2_buf_8 fanout2910 (.A(\data_pdata[19]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2910));
 sg13g2_buf_8 fanout2911 (.A(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2911));
 sg13g2_buf_8 fanout2912 (.A(\data_pdata[18]_sg13g2_mux2_1_A0_X_sg13g2_a21oi_1_A2_Y ),
    .X(net2912));
 sg13g2_buf_8 fanout2913 (.A(net2914),
    .X(net2913));
 sg13g2_buf_8 fanout2914 (.A(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y),
    .X(net2914));
 sg13g2_buf_8 fanout2915 (.A(net2917),
    .X(net2915));
 sg13g2_buf_1 fanout2916 (.A(net2917),
    .X(net2916));
 sg13g2_buf_8 fanout2917 (.A(target_sel_q_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_A_N_Y),
    .X(net2917));
 sg13g2_buf_8 fanout2918 (.A(net81),
    .X(net2918));
 sg13g2_buf_8 fanout2919 (.A(net81),
    .X(net2919));
 sg13g2_buf_16 fanout2920 (.X(net2920),
    .A(net2921));
 sg13g2_buf_8 fanout2921 (.A(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_A2 ),
    .X(net2921));
 sg13g2_buf_8 fanout2922 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D ),
    .X(net2922));
 sg13g2_buf_8 fanout2923 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand4_1_Y_C ),
    .X(net2923));
 sg13g2_buf_8 fanout2924 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2 ),
    .X(net2924));
 sg13g2_buf_8 fanout2925 (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q_sg13g2_a21oi_1_A1_A2_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B),
    .X(net2925));
 sg13g2_buf_8 fanout2926 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y ),
    .X(net2926));
 sg13g2_buf_8 fanout2927 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2927));
 sg13g2_buf_8 fanout2928 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2928));
 sg13g2_buf_8 fanout2929 (.A(net2932),
    .X(net2929));
 sg13g2_buf_8 fanout2930 (.A(net2932),
    .X(net2930));
 sg13g2_buf_8 fanout2931 (.A(net2932),
    .X(net2931));
 sg13g2_buf_8 fanout2932 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2932));
 sg13g2_buf_8 fanout2933 (.A(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2 ),
    .X(net2933));
 sg13g2_buf_8 fanout2934 (.A(\i_snitch.inst_addr_o[18]_sg13g2_a221oi_1_A1_B2_sg13g2_a221oi_1_Y_B2 ),
    .X(net2934));
 sg13g2_buf_8 fanout2935 (.A(net2939),
    .X(net2935));
 sg13g2_buf_8 fanout2936 (.A(net2938),
    .X(net2936));
 sg13g2_buf_8 fanout2937 (.A(net2938),
    .X(net2937));
 sg13g2_buf_8 fanout2938 (.A(net2939),
    .X(net2938));
 sg13g2_buf_8 fanout2939 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2939));
 sg13g2_buf_8 fanout2940 (.A(net2941),
    .X(net2940));
 sg13g2_buf_8 fanout2941 (.A(net2946),
    .X(net2941));
 sg13g2_buf_8 fanout2942 (.A(net2945),
    .X(net2942));
 sg13g2_buf_2 fanout2943 (.A(net2945),
    .X(net2943));
 sg13g2_buf_8 fanout2944 (.A(net2945),
    .X(net2944));
 sg13g2_buf_8 fanout2945 (.A(net2946),
    .X(net2945));
 sg13g2_buf_8 fanout2946 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net2946));
 sg13g2_buf_8 fanout2947 (.A(net2949),
    .X(net2947));
 sg13g2_buf_8 fanout2948 (.A(net2949),
    .X(net2948));
 sg13g2_buf_8 fanout2949 (.A(net111),
    .X(net2949));
 sg13g2_buf_8 fanout2950 (.A(net2951),
    .X(net2950));
 sg13g2_buf_8 fanout2951 (.A(net2953),
    .X(net2951));
 sg13g2_buf_8 fanout2952 (.A(net2953),
    .X(net2952));
 sg13g2_buf_8 fanout2953 (.A(net111),
    .X(net2953));
 sg13g2_buf_8 fanout2954 (.A(net2955),
    .X(net2954));
 sg13g2_buf_8 fanout2955 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net2955));
 sg13g2_buf_8 fanout2956 (.A(net2960),
    .X(net2956));
 sg13g2_buf_2 fanout2957 (.A(net2960),
    .X(net2957));
 sg13g2_buf_8 fanout2958 (.A(net2960),
    .X(net2958));
 sg13g2_buf_8 fanout2959 (.A(net2960),
    .X(net2959));
 sg13g2_buf_8 fanout2960 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2960));
 sg13g2_buf_8 fanout2961 (.A(net2962),
    .X(net2961));
 sg13g2_buf_8 fanout2962 (.A(net2967),
    .X(net2962));
 sg13g2_buf_8 fanout2963 (.A(net2966),
    .X(net2963));
 sg13g2_buf_8 fanout2964 (.A(net2966),
    .X(net2964));
 sg13g2_buf_8 fanout2965 (.A(net2966),
    .X(net2965));
 sg13g2_buf_8 fanout2966 (.A(net2967),
    .X(net2966));
 sg13g2_buf_8 fanout2967 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net2967));
 sg13g2_buf_8 fanout2968 (.A(net2969),
    .X(net2968));
 sg13g2_buf_8 fanout2969 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2969));
 sg13g2_buf_8 fanout2970 (.A(net2972),
    .X(net2970));
 sg13g2_buf_8 fanout2971 (.A(net2972),
    .X(net2971));
 sg13g2_buf_8 fanout2972 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2972));
 sg13g2_buf_8 fanout2973 (.A(net2976),
    .X(net2973));
 sg13g2_buf_8 fanout2974 (.A(net2976),
    .X(net2974));
 sg13g2_buf_1 fanout2975 (.A(net2976),
    .X(net2975));
 sg13g2_buf_8 fanout2976 (.A(net2996),
    .X(net2976));
 sg13g2_buf_8 fanout2977 (.A(net2979),
    .X(net2977));
 sg13g2_buf_8 fanout2978 (.A(net2979),
    .X(net2978));
 sg13g2_buf_8 fanout2979 (.A(net2996),
    .X(net2979));
 sg13g2_buf_8 fanout2980 (.A(net2984),
    .X(net2980));
 sg13g2_buf_1 fanout2981 (.A(net2984),
    .X(net2981));
 sg13g2_buf_8 fanout2982 (.A(net2984),
    .X(net2982));
 sg13g2_buf_8 fanout2983 (.A(net2984),
    .X(net2983));
 sg13g2_buf_8 fanout2984 (.A(net2996),
    .X(net2984));
 sg13g2_buf_8 fanout2985 (.A(net2986),
    .X(net2985));
 sg13g2_buf_8 fanout2986 (.A(net2995),
    .X(net2986));
 sg13g2_buf_8 fanout2987 (.A(net2989),
    .X(net2987));
 sg13g2_buf_8 fanout2988 (.A(net2989),
    .X(net2988));
 sg13g2_buf_8 fanout2989 (.A(net2995),
    .X(net2989));
 sg13g2_buf_8 fanout2990 (.A(net2995),
    .X(net2990));
 sg13g2_buf_8 fanout2991 (.A(net2995),
    .X(net2991));
 sg13g2_buf_8 fanout2992 (.A(net2994),
    .X(net2992));
 sg13g2_buf_8 fanout2993 (.A(net2994),
    .X(net2993));
 sg13g2_buf_8 fanout2994 (.A(net2995),
    .X(net2994));
 sg13g2_buf_8 fanout2995 (.A(net2996),
    .X(net2995));
 sg13g2_buf_8 fanout2996 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net2996));
 sg13g2_buf_8 fanout2997 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2997));
 sg13g2_buf_8 fanout2998 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net2998));
 sg13g2_buf_8 fanout2999 (.A(net3003),
    .X(net2999));
 sg13g2_buf_8 fanout3000 (.A(net3003),
    .X(net3000));
 sg13g2_buf_8 fanout3001 (.A(net3003),
    .X(net3001));
 sg13g2_buf_1 fanout3002 (.A(net3003),
    .X(net3002));
 sg13g2_buf_8 fanout3003 (.A(net3011),
    .X(net3003));
 sg13g2_buf_8 fanout3004 (.A(net3006),
    .X(net3004));
 sg13g2_buf_8 fanout3005 (.A(net3006),
    .X(net3005));
 sg13g2_buf_8 fanout3006 (.A(net3011),
    .X(net3006));
 sg13g2_buf_8 fanout3007 (.A(net3010),
    .X(net3007));
 sg13g2_buf_8 fanout3008 (.A(net3009),
    .X(net3008));
 sg13g2_buf_8 fanout3009 (.A(net3010),
    .X(net3009));
 sg13g2_buf_8 fanout3010 (.A(net3011),
    .X(net3010));
 sg13g2_buf_8 fanout3011 (.A(net3025),
    .X(net3011));
 sg13g2_buf_8 fanout3012 (.A(net3015),
    .X(net3012));
 sg13g2_buf_8 fanout3013 (.A(net3015),
    .X(net3013));
 sg13g2_buf_8 fanout3014 (.A(net3015),
    .X(net3014));
 sg13g2_buf_8 fanout3015 (.A(net3025),
    .X(net3015));
 sg13g2_buf_8 fanout3016 (.A(net3018),
    .X(net3016));
 sg13g2_buf_8 fanout3017 (.A(net3018),
    .X(net3017));
 sg13g2_buf_8 fanout3018 (.A(net3025),
    .X(net3018));
 sg13g2_buf_8 fanout3019 (.A(net3024),
    .X(net3019));
 sg13g2_buf_8 fanout3020 (.A(net3021),
    .X(net3020));
 sg13g2_buf_8 fanout3021 (.A(net3023),
    .X(net3021));
 sg13g2_buf_8 fanout3022 (.A(net3023),
    .X(net3022));
 sg13g2_buf_8 fanout3023 (.A(net3024),
    .X(net3023));
 sg13g2_buf_8 fanout3024 (.A(net3025),
    .X(net3024));
 sg13g2_buf_8 fanout3025 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nor2b_1_B_N_Y ),
    .X(net3025));
 sg13g2_buf_8 fanout3026 (.A(net3027),
    .X(net3026));
 sg13g2_buf_8 fanout3027 (.A(net3032),
    .X(net3027));
 sg13g2_buf_8 fanout3028 (.A(net3031),
    .X(net3028));
 sg13g2_buf_8 fanout3029 (.A(net3031),
    .X(net3029));
 sg13g2_buf_8 fanout3030 (.A(net3031),
    .X(net3030));
 sg13g2_buf_8 fanout3031 (.A(net3032),
    .X(net3031));
 sg13g2_buf_8 fanout3032 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_nand2b_1_A_N_Y_sg13g2_nand2b_1_B_Y ),
    .X(net3032));
 sg13g2_buf_8 fanout3033 (.A(net3034),
    .X(net3033));
 sg13g2_buf_8 fanout3034 (.A(net3037),
    .X(net3034));
 sg13g2_buf_2 fanout3035 (.A(net3037),
    .X(net3035));
 sg13g2_buf_1 fanout3036 (.A(net3037),
    .X(net3036));
 sg13g2_buf_2 fanout3037 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_1_Y ),
    .X(net3037));
 sg13g2_buf_8 fanout3038 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y),
    .X(net3038));
 sg13g2_buf_8 fanout3039 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y),
    .X(net3039));
 sg13g2_buf_8 fanout3040 (.A(net3042),
    .X(net3040));
 sg13g2_buf_8 fanout3041 (.A(net3042),
    .X(net3041));
 sg13g2_buf_8 fanout3042 (.A(data_pvalid_sg13g2_nand2b_1_B_Y_sg13g2_nor4_1_C_Y),
    .X(net3042));
 sg13g2_buf_8 fanout3043 (.A(net3044),
    .X(net3043));
 sg13g2_buf_8 fanout3044 (.A(net3045),
    .X(net3044));
 sg13g2_buf_8 fanout3045 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X ),
    .X(net3045));
 sg13g2_buf_8 fanout3046 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X ),
    .X(net3046));
 sg13g2_buf_2 fanout3047 (.A(\cnt_q[2]_sg13g2_nand3_1_A_Y_sg13g2_and2_1_B_X ),
    .X(net3047));
 sg13g2_buf_8 fanout3048 (.A(net3049),
    .X(net3048));
 sg13g2_buf_8 fanout3049 (.A(net3052),
    .X(net3049));
 sg13g2_buf_8 fanout3050 (.A(net3051),
    .X(net3050));
 sg13g2_buf_8 fanout3051 (.A(net3052),
    .X(net3051));
 sg13g2_buf_8 fanout3052 (.A(target_sel_q_sg13g2_nand2_1_B_Y),
    .X(net3052));
 sg13g2_buf_8 fanout3053 (.A(net3055),
    .X(net3053));
 sg13g2_buf_1 fanout3054 (.A(net3055),
    .X(net3054));
 sg13g2_buf_8 fanout3055 (.A(state_sg13g2_inv_1_A_Y),
    .X(net3055));
 sg13g2_buf_8 fanout3056 (.A(state_sg13g2_inv_1_A_Y),
    .X(net3056));
 sg13g2_buf_1 fanout3057 (.A(state_sg13g2_inv_1_A_Y),
    .X(net3057));
 sg13g2_buf_8 fanout3058 (.A(net3059),
    .X(net3058));
 sg13g2_buf_8 fanout3059 (.A(net3062),
    .X(net3059));
 sg13g2_buf_8 fanout3060 (.A(net3061),
    .X(net3060));
 sg13g2_buf_8 fanout3061 (.A(net3062),
    .X(net3061));
 sg13g2_buf_2 fanout3062 (.A(rsp_state_q_sg13g2_nor2_1_A_Y),
    .X(net3062));
 sg13g2_buf_8 fanout3063 (.A(net3064),
    .X(net3063));
 sg13g2_buf_8 fanout3064 (.A(net3067),
    .X(net3064));
 sg13g2_buf_8 fanout3065 (.A(net3067),
    .X(net3065));
 sg13g2_buf_8 fanout3066 (.A(net3067),
    .X(net3066));
 sg13g2_buf_8 fanout3067 (.A(rsp_data_ready),
    .X(net3067));
 sg13g2_buf_8 fanout3068 (.A(net3069),
    .X(net3068));
 sg13g2_buf_8 fanout3069 (.A(\i_snitch.i_snitch_lsu.metadata_q[1]_sg13g2_nand2b_1_B_Y ),
    .X(net3069));
 sg13g2_buf_8 fanout3070 (.A(\i_snitch.i_snitch_lsu.metadata_q[0]_sg13g2_or2_1_A_X ),
    .X(net3070));
 sg13g2_buf_8 fanout3071 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_mux2_1_A1_1_X ),
    .X(net3071));
 sg13g2_buf_8 fanout3072 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_mux2_1_A1_1_X ),
    .X(net3072));
 sg13g2_buf_8 fanout3073 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_mux2_1_A1_X ),
    .X(net3073));
 sg13g2_buf_8 fanout3074 (.A(net3075),
    .X(net3074));
 sg13g2_buf_8 fanout3075 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_mux2_1_A1_X ),
    .X(net3075));
 sg13g2_buf_8 fanout3076 (.A(net3077),
    .X(net3076));
 sg13g2_buf_8 fanout3077 (.A(net3078),
    .X(net3077));
 sg13g2_buf_8 fanout3078 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_mux2_1_A1_1_X ),
    .X(net3078));
 sg13g2_buf_8 fanout3079 (.A(net3080),
    .X(net3079));
 sg13g2_buf_8 fanout3080 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_mux2_1_A1_1_X ),
    .X(net3080));
 sg13g2_buf_8 fanout3081 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ),
    .X(net3081));
 sg13g2_buf_8 fanout3082 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_mux2_1_A1_1_X ),
    .X(net3082));
 sg13g2_buf_8 fanout3083 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_X ),
    .X(net3083));
 sg13g2_buf_1 fanout3084 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_mux2_1_A1_X ),
    .X(net3084));
 sg13g2_buf_8 fanout3085 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ),
    .X(net3085));
 sg13g2_buf_1 fanout3086 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_mux2_1_A1_1_X ),
    .X(net3086));
 sg13g2_buf_8 fanout3087 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_mux2_1_A1_1_X ),
    .X(net3087));
 sg13g2_buf_8 fanout3088 (.A(net3090),
    .X(net3088));
 sg13g2_buf_8 fanout3089 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_X ),
    .X(net3089));
 sg13g2_buf_8 fanout3090 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_mux2_1_A1_X ),
    .X(net3090));
 sg13g2_buf_8 fanout3091 (.A(net3093),
    .X(net3091));
 sg13g2_buf_2 fanout3092 (.A(net3093),
    .X(net3092));
 sg13g2_buf_8 fanout3093 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_X ),
    .X(net3093));
 sg13g2_buf_8 fanout3094 (.A(net3097),
    .X(net3094));
 sg13g2_buf_2 fanout3095 (.A(net3097),
    .X(net3095));
 sg13g2_buf_8 fanout3096 (.A(net3097),
    .X(net3096));
 sg13g2_buf_8 fanout3097 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_mux2_1_A1_X ),
    .X(net3097));
 sg13g2_buf_8 fanout3098 (.A(net3099),
    .X(net3098));
 sg13g2_buf_8 fanout3099 (.A(net3102),
    .X(net3099));
 sg13g2_buf_8 fanout3100 (.A(net3101),
    .X(net3100));
 sg13g2_buf_8 fanout3101 (.A(net3102),
    .X(net3101));
 sg13g2_buf_8 fanout3102 (.A(net3105),
    .X(net3102));
 sg13g2_buf_8 fanout3103 (.A(net3105),
    .X(net3103));
 sg13g2_buf_8 fanout3104 (.A(net3105),
    .X(net3104));
 sg13g2_buf_8 fanout3105 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_X ),
    .X(net3105));
 sg13g2_buf_8 fanout3106 (.A(net3107),
    .X(net3106));
 sg13g2_buf_8 fanout3107 (.A(net3110),
    .X(net3107));
 sg13g2_buf_8 fanout3108 (.A(net3110),
    .X(net3108));
 sg13g2_buf_8 fanout3109 (.A(net3110),
    .X(net3109));
 sg13g2_buf_8 fanout3110 (.A(net3114),
    .X(net3110));
 sg13g2_buf_8 fanout3111 (.A(net3114),
    .X(net3111));
 sg13g2_buf_8 fanout3112 (.A(net3114),
    .X(net3112));
 sg13g2_buf_8 fanout3113 (.A(net3114),
    .X(net3113));
 sg13g2_buf_16 fanout3114 (.X(net3114),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_mux2_1_A1_X ));
 sg13g2_buf_8 fanout3115 (.A(net3118),
    .X(net3115));
 sg13g2_buf_8 fanout3116 (.A(net3118),
    .X(net3116));
 sg13g2_buf_8 fanout3117 (.A(net3118),
    .X(net3117));
 sg13g2_buf_8 fanout3118 (.A(net3121),
    .X(net3118));
 sg13g2_buf_8 fanout3119 (.A(net3120),
    .X(net3119));
 sg13g2_buf_8 fanout3120 (.A(net3121),
    .X(net3120));
 sg13g2_buf_8 fanout3121 (.A(net79),
    .X(net3121));
 sg13g2_buf_8 fanout3122 (.A(net3125),
    .X(net3122));
 sg13g2_buf_8 fanout3123 (.A(net3125),
    .X(net3123));
 sg13g2_buf_8 fanout3124 (.A(net3125),
    .X(net3124));
 sg13g2_buf_8 fanout3125 (.A(net80),
    .X(net3125));
 sg13g2_buf_8 fanout3126 (.A(net3128),
    .X(net3126));
 sg13g2_buf_8 fanout3127 (.A(net3128),
    .X(net3127));
 sg13g2_buf_16 fanout3128 (.X(net3128),
    .A(net3132));
 sg13g2_buf_8 fanout3129 (.A(net3131),
    .X(net3129));
 sg13g2_buf_8 fanout3130 (.A(net3131),
    .X(net3130));
 sg13g2_buf_8 fanout3131 (.A(net3132),
    .X(net3131));
 sg13g2_buf_16 fanout3132 (.X(net3132),
    .A(net3140));
 sg13g2_buf_8 fanout3133 (.A(net107),
    .X(net3133));
 sg13g2_buf_8 fanout3134 (.A(net3140),
    .X(net3134));
 sg13g2_buf_8 fanout3135 (.A(net3139),
    .X(net3135));
 sg13g2_buf_8 fanout3136 (.A(net3139),
    .X(net3136));
 sg13g2_buf_8 fanout3137 (.A(net3139),
    .X(net3137));
 sg13g2_buf_8 fanout3138 (.A(net3139),
    .X(net3138));
 sg13g2_buf_8 fanout3139 (.A(net3140),
    .X(net3139));
 sg13g2_buf_16 fanout3140 (.X(net3140),
    .A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_X ));
 sg13g2_buf_8 fanout3141 (.A(net109),
    .X(net3141));
 sg13g2_buf_8 fanout3142 (.A(net3143),
    .X(net3142));
 sg13g2_buf_8 fanout3143 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ),
    .X(net3143));
 sg13g2_buf_8 fanout3144 (.A(net3146),
    .X(net3144));
 sg13g2_buf_8 fanout3145 (.A(net3146),
    .X(net3145));
 sg13g2_buf_8 fanout3146 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_X ),
    .X(net3146));
 sg13g2_buf_8 fanout3147 (.A(net3148),
    .X(net3147));
 sg13g2_buf_8 fanout3148 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_mux2_1_A1_X ),
    .X(net3148));
 sg13g2_buf_8 fanout3149 (.A(net3150),
    .X(net3149));
 sg13g2_buf_8 fanout3150 (.A(net3151),
    .X(net3150));
 sg13g2_buf_8 fanout3151 (.A(\i_snitch.i_snitch_lsu.metadata_q[3] ),
    .X(net3151));
 sg13g2_buf_8 fanout3152 (.A(net3153),
    .X(net3152));
 sg13g2_buf_8 fanout3153 (.A(net3154),
    .X(net3153));
 sg13g2_buf_8 fanout3154 (.A(net1403),
    .X(net3154));
 sg13g2_buf_8 fanout3155 (.A(net3158),
    .X(net3155));
 sg13g2_buf_1 fanout3156 (.A(net3157),
    .X(net3156));
 sg13g2_buf_2 fanout3157 (.A(net3158),
    .X(net3157));
 sg13g2_buf_8 fanout3158 (.A(\i_snitch.i_snitch_lsu.metadata_q[2] ),
    .X(net3158));
 sg13g2_buf_2 fanout3159 (.A(net3160),
    .X(net3159));
 sg13g2_buf_2 fanout3160 (.A(net3161),
    .X(net3160));
 sg13g2_buf_1 fanout3161 (.A(net3162),
    .X(net3161));
 sg13g2_buf_8 fanout3162 (.A(net1404),
    .X(net3162));
 sg13g2_buf_8 fanout3163 (.A(net1402),
    .X(net3163));
 sg13g2_buf_8 fanout3164 (.A(net3165),
    .X(net3164));
 sg13g2_buf_8 fanout3165 (.A(net3167),
    .X(net3165));
 sg13g2_buf_8 fanout3166 (.A(net3167),
    .X(net3166));
 sg13g2_buf_8 fanout3167 (.A(net3173),
    .X(net3167));
 sg13g2_buf_8 fanout3168 (.A(net3173),
    .X(net3168));
 sg13g2_buf_8 fanout3169 (.A(net3171),
    .X(net3169));
 sg13g2_buf_8 fanout3170 (.A(net3171),
    .X(net3170));
 sg13g2_buf_8 fanout3171 (.A(net3172),
    .X(net3171));
 sg13g2_buf_8 fanout3172 (.A(net3173),
    .X(net3172));
 sg13g2_buf_8 fanout3173 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_full_q ),
    .X(net3173));
 sg13g2_buf_8 fanout3174 (.A(net3176),
    .X(net3174));
 sg13g2_buf_8 fanout3175 (.A(net3176),
    .X(net3175));
 sg13g2_buf_16 fanout3176 (.X(net3176),
    .A(net3183));
 sg13g2_buf_8 fanout3177 (.A(net105),
    .X(net3177));
 sg13g2_buf_8 fanout3178 (.A(net3182),
    .X(net3178));
 sg13g2_buf_8 fanout3179 (.A(net3180),
    .X(net3179));
 sg13g2_buf_16 fanout3180 (.X(net3180),
    .A(net3181));
 sg13g2_buf_16 fanout3181 (.X(net3181),
    .A(net3182));
 sg13g2_buf_16 fanout3182 (.X(net3182),
    .A(net3183));
 sg13g2_buf_8 fanout3183 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q ),
    .X(net3183));
 sg13g2_buf_8 fanout3184 (.A(net3194),
    .X(net3184));
 sg13g2_buf_8 fanout3185 (.A(net3194),
    .X(net3185));
 sg13g2_buf_8 fanout3186 (.A(net3188),
    .X(net3186));
 sg13g2_buf_8 fanout3187 (.A(net3188),
    .X(net3187));
 sg13g2_buf_8 fanout3188 (.A(net3194),
    .X(net3188));
 sg13g2_buf_8 fanout3189 (.A(net3193),
    .X(net3189));
 sg13g2_buf_8 fanout3190 (.A(net3193),
    .X(net3190));
 sg13g2_buf_8 fanout3191 (.A(net3193),
    .X(net3191));
 sg13g2_buf_8 fanout3192 (.A(net3193),
    .X(net3192));
 sg13g2_buf_8 fanout3193 (.A(net3194),
    .X(net3193));
 sg13g2_buf_8 fanout3194 (.A(net3226),
    .X(net3194));
 sg13g2_buf_8 fanout3195 (.A(net3197),
    .X(net3195));
 sg13g2_buf_8 fanout3196 (.A(net3197),
    .X(net3196));
 sg13g2_buf_8 fanout3197 (.A(net3205),
    .X(net3197));
 sg13g2_buf_8 fanout3198 (.A(net3200),
    .X(net3198));
 sg13g2_buf_8 fanout3199 (.A(net3200),
    .X(net3199));
 sg13g2_buf_8 fanout3200 (.A(net3205),
    .X(net3200));
 sg13g2_buf_8 fanout3201 (.A(net3202),
    .X(net3201));
 sg13g2_buf_8 fanout3202 (.A(net3205),
    .X(net3202));
 sg13g2_buf_8 fanout3203 (.A(net3205),
    .X(net3203));
 sg13g2_buf_2 fanout3204 (.A(net3205),
    .X(net3204));
 sg13g2_buf_8 fanout3205 (.A(net3226),
    .X(net3205));
 sg13g2_buf_8 fanout3206 (.A(net3208),
    .X(net3206));
 sg13g2_buf_8 fanout3207 (.A(net3211),
    .X(net3207));
 sg13g2_buf_2 fanout3208 (.A(net3211),
    .X(net3208));
 sg13g2_buf_8 fanout3209 (.A(net3210),
    .X(net3209));
 sg13g2_buf_8 fanout3210 (.A(net3211),
    .X(net3210));
 sg13g2_buf_8 fanout3211 (.A(net3226),
    .X(net3211));
 sg13g2_buf_8 fanout3212 (.A(net3213),
    .X(net3212));
 sg13g2_buf_8 fanout3213 (.A(net3216),
    .X(net3213));
 sg13g2_buf_8 fanout3214 (.A(net3216),
    .X(net3214));
 sg13g2_buf_8 fanout3215 (.A(net3216),
    .X(net3215));
 sg13g2_buf_8 fanout3216 (.A(net3226),
    .X(net3216));
 sg13g2_buf_8 fanout3217 (.A(net3225),
    .X(net3217));
 sg13g2_buf_8 fanout3218 (.A(net3225),
    .X(net3218));
 sg13g2_buf_8 fanout3219 (.A(net3220),
    .X(net3219));
 sg13g2_buf_8 fanout3220 (.A(net3225),
    .X(net3220));
 sg13g2_buf_8 fanout3221 (.A(net3222),
    .X(net3221));
 sg13g2_buf_8 fanout3222 (.A(net3224),
    .X(net3222));
 sg13g2_buf_8 fanout3223 (.A(net3224),
    .X(net3223));
 sg13g2_buf_8 fanout3224 (.A(net3225),
    .X(net3224));
 sg13g2_buf_8 fanout3225 (.A(net3226),
    .X(net3225));
 sg13g2_buf_8 fanout3226 (.A(net3330),
    .X(net3226));
 sg13g2_buf_8 fanout3227 (.A(net3229),
    .X(net3227));
 sg13g2_buf_8 fanout3228 (.A(net3229),
    .X(net3228));
 sg13g2_buf_8 fanout3229 (.A(net3249),
    .X(net3229));
 sg13g2_buf_8 fanout3230 (.A(net3232),
    .X(net3230));
 sg13g2_buf_8 fanout3231 (.A(net3232),
    .X(net3231));
 sg13g2_buf_8 fanout3232 (.A(net3249),
    .X(net3232));
 sg13g2_buf_8 fanout3233 (.A(net3236),
    .X(net3233));
 sg13g2_buf_8 fanout3234 (.A(net3236),
    .X(net3234));
 sg13g2_buf_8 fanout3235 (.A(net3236),
    .X(net3235));
 sg13g2_buf_8 fanout3236 (.A(net3249),
    .X(net3236));
 sg13g2_buf_8 fanout3237 (.A(net3239),
    .X(net3237));
 sg13g2_buf_8 fanout3238 (.A(net3239),
    .X(net3238));
 sg13g2_buf_8 fanout3239 (.A(net3249),
    .X(net3239));
 sg13g2_buf_8 fanout3240 (.A(net3241),
    .X(net3240));
 sg13g2_buf_8 fanout3241 (.A(net3249),
    .X(net3241));
 sg13g2_buf_8 fanout3242 (.A(net3243),
    .X(net3242));
 sg13g2_buf_8 fanout3243 (.A(net3248),
    .X(net3243));
 sg13g2_buf_8 fanout3244 (.A(net3247),
    .X(net3244));
 sg13g2_buf_8 fanout3245 (.A(net3247),
    .X(net3245));
 sg13g2_buf_8 fanout3246 (.A(net3247),
    .X(net3246));
 sg13g2_buf_8 fanout3247 (.A(net3248),
    .X(net3247));
 sg13g2_buf_8 fanout3248 (.A(net3249),
    .X(net3248));
 sg13g2_buf_8 fanout3249 (.A(net3330),
    .X(net3249));
 sg13g2_buf_8 fanout3250 (.A(net3259),
    .X(net3250));
 sg13g2_buf_8 fanout3251 (.A(net3259),
    .X(net3251));
 sg13g2_buf_8 fanout3252 (.A(net3253),
    .X(net3252));
 sg13g2_buf_8 fanout3253 (.A(net3259),
    .X(net3253));
 sg13g2_buf_8 fanout3254 (.A(net3258),
    .X(net3254));
 sg13g2_buf_8 fanout3255 (.A(net3258),
    .X(net3255));
 sg13g2_buf_8 fanout3256 (.A(net3258),
    .X(net3256));
 sg13g2_buf_2 fanout3257 (.A(net3258),
    .X(net3257));
 sg13g2_buf_8 fanout3258 (.A(net3259),
    .X(net3258));
 sg13g2_buf_8 fanout3259 (.A(net3261),
    .X(net3259));
 sg13g2_buf_8 fanout3260 (.A(net3261),
    .X(net3260));
 sg13g2_buf_8 fanout3261 (.A(net3330),
    .X(net3261));
 sg13g2_buf_8 fanout3262 (.A(net3264),
    .X(net3262));
 sg13g2_buf_8 fanout3263 (.A(net3264),
    .X(net3263));
 sg13g2_buf_8 fanout3264 (.A(net3272),
    .X(net3264));
 sg13g2_buf_8 fanout3265 (.A(net3272),
    .X(net3265));
 sg13g2_buf_8 fanout3266 (.A(net3272),
    .X(net3266));
 sg13g2_buf_8 fanout3267 (.A(net3268),
    .X(net3267));
 sg13g2_buf_8 fanout3268 (.A(net3271),
    .X(net3268));
 sg13g2_buf_8 fanout3269 (.A(net3271),
    .X(net3269));
 sg13g2_buf_8 fanout3270 (.A(net3271),
    .X(net3270));
 sg13g2_buf_8 fanout3271 (.A(net3272),
    .X(net3271));
 sg13g2_buf_8 fanout3272 (.A(net3329),
    .X(net3272));
 sg13g2_buf_8 fanout3273 (.A(net3282),
    .X(net3273));
 sg13g2_buf_8 fanout3274 (.A(net3282),
    .X(net3274));
 sg13g2_buf_8 fanout3275 (.A(net3276),
    .X(net3275));
 sg13g2_buf_8 fanout3276 (.A(net3282),
    .X(net3276));
 sg13g2_buf_8 fanout3277 (.A(net3281),
    .X(net3277));
 sg13g2_buf_8 fanout3278 (.A(net3281),
    .X(net3278));
 sg13g2_buf_8 fanout3279 (.A(net3281),
    .X(net3279));
 sg13g2_buf_8 fanout3280 (.A(net3281),
    .X(net3280));
 sg13g2_buf_8 fanout3281 (.A(net3282),
    .X(net3281));
 sg13g2_buf_8 fanout3282 (.A(net3329),
    .X(net3282));
 sg13g2_buf_8 fanout3283 (.A(net3284),
    .X(net3283));
 sg13g2_buf_8 fanout3284 (.A(net3287),
    .X(net3284));
 sg13g2_buf_8 fanout3285 (.A(net3287),
    .X(net3285));
 sg13g2_buf_8 fanout3286 (.A(net3287),
    .X(net3286));
 sg13g2_buf_8 fanout3287 (.A(net3301),
    .X(net3287));
 sg13g2_buf_8 fanout3288 (.A(net3301),
    .X(net3288));
 sg13g2_buf_8 fanout3289 (.A(net3290),
    .X(net3289));
 sg13g2_buf_8 fanout3290 (.A(net3301),
    .X(net3290));
 sg13g2_buf_8 fanout3291 (.A(net3300),
    .X(net3291));
 sg13g2_buf_8 fanout3292 (.A(net3300),
    .X(net3292));
 sg13g2_buf_8 fanout3293 (.A(net3294),
    .X(net3293));
 sg13g2_buf_8 fanout3294 (.A(net3300),
    .X(net3294));
 sg13g2_buf_8 fanout3295 (.A(net3300),
    .X(net3295));
 sg13g2_buf_8 fanout3296 (.A(net3300),
    .X(net3296));
 sg13g2_buf_8 fanout3297 (.A(net3299),
    .X(net3297));
 sg13g2_buf_8 fanout3298 (.A(net3299),
    .X(net3298));
 sg13g2_buf_8 fanout3299 (.A(net3300),
    .X(net3299));
 sg13g2_buf_8 fanout3300 (.A(net3301),
    .X(net3300));
 sg13g2_buf_8 fanout3301 (.A(net3329),
    .X(net3301));
 sg13g2_buf_8 fanout3302 (.A(net3306),
    .X(net3302));
 sg13g2_buf_8 fanout3303 (.A(net3306),
    .X(net3303));
 sg13g2_buf_8 fanout3304 (.A(net3306),
    .X(net3304));
 sg13g2_buf_8 fanout3305 (.A(net3306),
    .X(net3305));
 sg13g2_buf_8 fanout3306 (.A(net3313),
    .X(net3306));
 sg13g2_buf_8 fanout3307 (.A(net3311),
    .X(net3307));
 sg13g2_buf_8 fanout3308 (.A(net3311),
    .X(net3308));
 sg13g2_buf_8 fanout3309 (.A(net3311),
    .X(net3309));
 sg13g2_buf_8 fanout3310 (.A(net3311),
    .X(net3310));
 sg13g2_buf_8 fanout3311 (.A(net3313),
    .X(net3311));
 sg13g2_buf_8 fanout3312 (.A(net3313),
    .X(net3312));
 sg13g2_buf_8 fanout3313 (.A(net3329),
    .X(net3313));
 sg13g2_buf_8 fanout3314 (.A(net3316),
    .X(net3314));
 sg13g2_buf_1 fanout3315 (.A(net3316),
    .X(net3315));
 sg13g2_buf_8 fanout3316 (.A(net3326),
    .X(net3316));
 sg13g2_buf_8 fanout3317 (.A(net3326),
    .X(net3317));
 sg13g2_buf_8 fanout3318 (.A(net3326),
    .X(net3318));
 sg13g2_buf_8 fanout3319 (.A(net3325),
    .X(net3319));
 sg13g2_buf_1 fanout3320 (.A(net3325),
    .X(net3320));
 sg13g2_buf_8 fanout3321 (.A(net3325),
    .X(net3321));
 sg13g2_buf_8 fanout3322 (.A(net3324),
    .X(net3322));
 sg13g2_buf_2 fanout3323 (.A(net3324),
    .X(net3323));
 sg13g2_buf_8 fanout3324 (.A(net3325),
    .X(net3324));
 sg13g2_buf_8 fanout3325 (.A(net3326),
    .X(net3325));
 sg13g2_buf_8 fanout3326 (.A(net3329),
    .X(net3326));
 sg13g2_buf_8 fanout3327 (.A(net3328),
    .X(net3327));
 sg13g2_buf_8 fanout3328 (.A(net3329),
    .X(net3328));
 sg13g2_buf_8 fanout3329 (.A(net3330),
    .X(net3329));
 sg13g2_buf_8 fanout3330 (.A(rst_n),
    .X(net3330));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[7]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_tiehi heichips25_snitch_wrapper_25 (.L_HI(net25));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_leaf_5_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_10_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_leaf_11_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_12_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_4_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_120_clk));
 sg13g2_inv_2 clkload12 (.A(clknet_leaf_110_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_19_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_16_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_leaf_107_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_27_clk));
 sg13g2_inv_1 clkload19 (.A(clknet_leaf_30_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_leaf_38_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_leaf_34_clk));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_18_clk));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_23_clk));
 sg13g2_inv_1 clkload24 (.A(clknet_leaf_17_clk));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_47_clk));
 sg13g2_inv_1 clkload26 (.A(clknet_leaf_48_clk));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_21_clk));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_22_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_31_clk));
 sg13g2_buf_8 clkload30 (.A(clknet_leaf_44_clk));
 sg13g2_inv_4 clkload31 (.A(clknet_leaf_45_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_leaf_98_clk));
 sg13g2_inv_1 clkload33 (.A(clknet_leaf_113_clk));
 sg13g2_buf_8 clkload34 (.A(clknet_leaf_100_clk));
 sg13g2_inv_4 clkload35 (.A(clknet_leaf_104_clk));
 sg13g2_inv_2 clkload36 (.A(clknet_leaf_105_clk));
 sg13g2_buf_8 clkload37 (.A(clknet_leaf_75_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_leaf_103_clk));
 sg13g2_inv_2 clkload39 (.A(clknet_leaf_92_clk));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_94_clk));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_87_clk));
 sg13g2_inv_2 clkload42 (.A(clknet_leaf_89_clk));
 sg13g2_inv_2 clkload43 (.A(clknet_leaf_90_clk));
 sg13g2_buf_8 clkload44 (.A(clknet_leaf_76_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_leaf_77_clk));
 sg13g2_inv_1 clkload46 (.A(clknet_leaf_78_clk));
 sg13g2_inv_4 clkload47 (.A(clknet_leaf_83_clk));
 sg13g2_inv_1 clkload48 (.A(clknet_leaf_50_clk));
 sg13g2_inv_2 clkload49 (.A(clknet_leaf_71_clk));
 sg13g2_buf_8 clkload50 (.A(clknet_leaf_106_clk));
 sg13g2_inv_1 clkload51 (.A(clknet_leaf_73_clk));
 sg13g2_buf_8 clkload52 (.A(clknet_leaf_74_clk));
 sg13g2_buf_8 clkload53 (.A(clknet_leaf_52_clk));
 sg13g2_inv_2 clkload54 (.A(clknet_leaf_53_clk));
 sg13g2_inv_1 clkload55 (.A(clknet_leaf_54_clk));
 sg13g2_inv_2 clkload56 (.A(clknet_leaf_66_clk));
 sg13g2_inv_1 clkload57 (.A(clknet_leaf_68_clk));
 sg13g2_inv_1 clkload58 (.A(clknet_leaf_64_clk));
 sg13g2_buf_8 clkload59 (.A(clknet_leaf_80_clk));
 sg13g2_inv_1 clkload60 (.A(clknet_leaf_81_clk));
 sg13g2_inv_1 clkload61 (.A(clknet_leaf_61_clk));
 sg13g2_inv_1 clkload62 (.A(clknet_leaf_62_clk));
 sg13g2_inv_2 clkload63 (.A(clknet_leaf_82_clk));
 sg13g2_inv_8 clkload64 (.A(clknet_leaf_55_clk));
 sg13g2_inv_2 clkload65 (.A(clknet_leaf_67_clk));
 sg13g2_inv_2 clkload66 (.A(clknet_leaf_56_clk));
 sg13g2_inv_2 clkload67 (.A(clknet_leaf_59_clk));
 sg13g2_buf_8 rebuffer1 (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_nand4_1_D_Y ),
    .X(net33));
 sg13g2_buf_2 rebuffer2 (.A(net33),
    .X(net34));
 sg13g2_buf_8 rebuffer3 (.A(\i_snitch.i_snitch_regfile.mem[65]_sg13g2_nor2_1_A_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a221oi_1_B1_Y ),
    .X(net35));
 sg13g2_buf_1 rebuffer4 (.A(net35),
    .X(net36));
 sg13g2_buf_1 rebuffer5 (.A(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ),
    .X(net37));
 sg13g2_buf_1 rebuffer6 (.A(\i_snitch.i_snitch_regfile.mem[265]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_a21oi_1_B1_Y_sg13g2_a221oi_1_C1_Y ),
    .X(net38));
 sg13g2_buf_2 rebuffer7 (.A(\i_snitch.i_snitch_regfile.mem[47]_sg13g2_a21oi_1_A1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_a22oi_1_B2_Y_sg13g2_and2_1_B_X_sg13g2_nand4_1_D_Y_sg13g2_nand2_1_B_Y_sg13g2_nand4_1_C_Y ),
    .X(net39));
 sg13g2_buf_8 rebuffer8 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_Y ),
    .X(net40));
 sg13g2_buf_8 rebuffer9 (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_nor3_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .X(net41));
 sg13g2_buf_1 rebuffer10 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y_sg13g2_a221oi_1_B2_Y_sg13g2_o21ai_1_A2_Y ),
    .X(net42));
 sg13g2_buf_1 rebuffer11 (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_nand4_1_A_Y_sg13g2_or4_1_D_X_sg13g2_or4_1_D_X_sg13g2_nand4_1_D_Y ),
    .X(net43));
 sg13g2_buf_2 rebuffer12 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_C1_Y ),
    .X(net44));
 sg13g2_buf_8 rebuffer13 (.A(\i_snitch.pc_d[4]_sg13g2_inv_1_Y_A_sg13g2_a21oi_1_Y_B1_sg13g2_nor3_1_Y_C_sg13g2_a22oi_1_Y_B1_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .X(net45));
 sg13g2_buf_2 rebuffer14 (.A(\i_snitch.pc_d[14]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_o21ai_1_Y_A2_sg13g2_nand4_1_B_D_sg13g2_nand2_1_Y_B_sg13g2_nand3b_1_Y_B ),
    .X(net46));
 sg13g2_buf_8 rebuffer15 (.A(\i_snitch.i_snitch_regfile.mem[130]_sg13g2_mux4_1_A0_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor3_1_C_Y_sg13g2_a221oi_1_C1_Y ),
    .X(net47));
 sg13g2_buf_2 rebuffer16 (.A(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y_sg13g2_nand4_1_A_Y ),
    .X(net48));
 sg13g2_buf_1 rebuffer17 (.A(\i_snitch.pc_d[0]_sg13g2_nand2_1_Y_B_sg13g2_nand3_1_Y_B ),
    .X(net49));
 sg13g2_buf_1 rebuffer18 (.A(\i_snitch.pc_d[18]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_a21oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .X(net50));
 sg13g2_buf_2 rebuffer19 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .X(net51));
 sg13g2_buf_1 rebuffer20 (.A(net51),
    .X(net52));
 sg13g2_buf_1 rebuffer21 (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A_sg13g2_xnor2_1_Y_B ),
    .X(net53));
 sg13g2_buf_1 rebuffer22 (.A(\i_snitch.pc_d[30]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2 ),
    .X(net54));
 sg13g2_buf_2 rebuffer23 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A_sg13g2_xor2_1_X_B_sg13g2_xor2_1_X_B ),
    .X(net55));
 sg13g2_buf_1 rebuffer24 (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1 ),
    .X(net56));
 sg13g2_buf_1 rebuffer25 (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1 ),
    .X(net57));
 sg13g2_buf_1 rebuffer26 (.A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand2_1_Y_A_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(net58));
 sg13g2_buf_1 rebuffer27 (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .X(net59));
 sg13g2_buf_1 rebuffer28 (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .X(net60));
 sg13g2_buf_1 rebuffer29 (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_mux4_1_A0_X_sg13g2_a21oi_1_A2_Y_sg13g2_a21o_1_A2_X_sg13g2_o21ai_1_A2_Y_sg13g2_nor2_1_B_Y_sg13g2_and4_1_D_A ),
    .X(net61));
 sg13g2_buf_1 rebuffer30 (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1 ),
    .X(net62));
 sg13g2_buf_1 rebuffer31 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net63));
 sg13g2_buf_1 rebuffer32 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_A1_sg13g2_xnor2_1_A_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net64));
 sg13g2_buf_1 rebuffer33 (.A(\i_snitch.i_snitch_regfile.mem[32]_sg13g2_a221oi_1_A1_Y_sg13g2_or2_1_A_X_sg13g2_a221oi_1_C1_Y_sg13g2_nor2b_1_A_Y ),
    .X(net65));
 sg13g2_buf_1 rebuffer34 (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nand4_1_Y_D_sg13g2_a22oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(net66));
 sg13g2_buf_1 rebuffer35 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_inv_1_Y_A ),
    .X(net67));
 sg13g2_buf_16 rebuffer36 (.X(net68),
    .A(net2241));
 sg13g2_buf_1 rebuffer37 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .X(net69));
 sg13g2_buf_2 rebuffer38 (.A(net40),
    .X(net70));
 sg13g2_buf_1 rebuffer39 (.A(\i_snitch.pc_d[19]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2 ),
    .X(net71));
 sg13g2_buf_1 rebuffer40 (.A(\i_snitch.pc_d[27]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_B ),
    .X(net72));
 sg13g2_buf_1 rebuffer41 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_mux2_1_A1_X ),
    .X(net73));
 sg13g2_buf_1 rebuffer42 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_mux2_1_A1_1_X ),
    .X(net74));
 sg13g2_buf_1 rebuffer43 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_A_sg13g2_nand3_1_B_Y_sg13g2_nor4_1_A_C_sg13g2_or2_1_B_A_sg13g2_a21o_1_B1_A2_sg13g2_a22oi_1_B1_Y ),
    .X(net75));
 sg13g2_buf_1 rebuffer44 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ),
    .X(net76));
 sg13g2_buf_1 rebuffer45 (.A(\i_snitch.pc_d[31]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a22oi_1_Y_A2_sg13g2_inv_1_Y_A ),
    .X(net77));
 sg13g2_buf_1 rebuffer46 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B_sg13g2_nand3_1_Y_B ),
    .X(net78));
 sg13g2_buf_1 rebuffer47 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_X ),
    .X(net79));
 sg13g2_buf_1 rebuffer48 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_mux2_1_A1_X ),
    .X(net80));
 sg13g2_buf_8 rebuffer49 (.A(\i_snitch.i_snitch_regfile.mem[129]_sg13g2_a22oi_1_A1_A2 ),
    .X(net81));
 sg13g2_buf_1 rebuffer50 (.A(\i_snitch.pc_d[3]_sg13g2_a21o_1_X_B1_sg13g2_and2_1_X_B_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .X(net82));
 sg13g2_buf_1 rebuffer51 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A1_sg13g2_nor2_1_Y_A ),
    .X(net83));
 sg13g2_buf_1 rebuffer52 (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .X(net84));
 sg13g2_buf_1 rebuffer53 (.A(\i_snitch.pc_d[15]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_A ),
    .X(net85));
 sg13g2_buf_1 rebuffer54 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_a221oi_1_A1_Y ),
    .X(net86));
 sg13g2_buf_1 rebuffer55 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_B1_sg13g2_nor4_1_Y_D_sg13g2_nor3_1_C_Y ),
    .X(net87));
 sg13g2_buf_1 rebuffer56 (.A(net2563),
    .X(net88));
 sg13g2_buf_1 rebuffer57 (.A(net2609),
    .X(net89));
 sg13g2_buf_1 rebuffer58 (.A(\i_snitch.i_snitch_regfile.mem[427]_sg13g2_inv_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_o21ai_1_A1_Y_sg13g2_o21ai_1_A2_Y_sg13g2_a21oi_1_B1_Y ),
    .X(net90));
 sg13g2_buf_1 rebuffer59 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_o21ai_1_B1_Y ),
    .X(net91));
 sg13g2_buf_1 rebuffer60 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_or3_1_C_X_sg13g2_a21o_1_B1_X ),
    .X(net92));
 sg13g2_buf_1 rebuffer61 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_a221oi_1_Y_B2 ),
    .X(net93));
 sg13g2_buf_1 rebuffer62 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y ),
    .X(net94));
 sg13g2_buf_2 rebuffer63 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_o21ai_1_B1_Y ),
    .X(net95));
 sg13g2_buf_2 rebuffer64 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_nand2_1_B_Y_sg13g2_and2_1_A_X_sg13g2_a221oi_1_B2_C1_sg13g2_nor3_1_Y_A ),
    .X(net96));
 sg13g2_buf_1 rebuffer65 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_nand3_1_A_Y_sg13g2_a221oi_1_A1_Y_sg13g2_and3_1_C_X_sg13g2_or2_1_B_X ),
    .X(net97));
 sg13g2_buf_1 rebuffer66 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_B_sg13g2_nor4_1_Y_C_sg13g2_a21o_1_X_A2_sg13g2_nor2b_1_Y_B_N_sg13g2_nand4_1_D_C_sg13g2_and4_1_X_C ),
    .X(net98));
 sg13g2_buf_1 rebuffer67 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_B ),
    .X(net99));
 sg13g2_buf_1 rebuffer68 (.A(net2537),
    .X(net100));
 sg13g2_buf_1 rebuffer69 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A ),
    .X(net101));
 sg13g2_buf_1 rebuffer70 (.A(\i_snitch.pc_d[12]_sg13g2_a22oi_1_Y_B2_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_a221oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_and4_1_D_C ),
    .X(net102));
 sg13g2_buf_1 rebuffer71 (.A(\i_snitch.pc_d[25]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_nor2_1_Y_B_sg13g2_nor2_1_Y_B_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B_sg13g2_xnor2_1_Y_A ),
    .X(net103));
 sg13g2_buf_1 rebuffer72 (.A(\i_snitch.pc_d[29]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_B1_sg13g2_a21oi_1_Y_A2_sg13g2_xor2_1_X_A_sg13g2_xor2_1_X_B ),
    .X(net104));
 sg13g2_buf_1 rebuffer73 (.A(net3183),
    .X(net105));
 sg13g2_buf_8 rebuffer74 (.A(net2311),
    .X(net106));
 sg13g2_buf_1 rebuffer75 (.A(net3140),
    .X(net107));
 sg13g2_buf_1 rebuffer76 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_mux2_1_A1_1_X_sg13g2_nor2b_1_A_Y ),
    .X(net108));
 sg13g2_buf_1 rebuffer77 (.A(net3143),
    .X(net109));
 sg13g2_buf_1 rebuffer78 (.A(net2921),
    .X(net110));
 sg13g2_buf_2 rebuffer79 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_nand2b_1_A_N_Y_sg13g2_o21ai_1_B1_Y ),
    .X(net111));
 sg13g2_buf_1 rebuffer80 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A2_sg13g2_nand4_1_Y_A_sg13g2_and4_1_A_X ),
    .X(net112));
 sg13g2_buf_1 rebuffer81 (.A(\i_snitch.i_snitch_regfile.mem[34]_sg13g2_a221oi_1_A1_Y_sg13g2_nor3_1_B_Y_sg13g2_o21ai_1_B1_A1_sg13g2_nand2_1_Y_A_sg13g2_and2_1_A_X ),
    .X(net113));
 sg13g2_buf_1 rebuffer82 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_mux2_1_A1_X ),
    .X(net114));
 sg13g2_buf_1 rebuffer83 (.A(\i_snitch.pc_d[2]_sg13g2_mux2_1_X_A1_sg13g2_o21ai_1_Y_B1_sg13g2_nand2_1_Y_B_sg13g2_a22oi_1_Y_A2_sg13g2_xnor2_1_Y_A_sg13g2_o21ai_1_A1_Y ),
    .X(net115));
 sg13g2_buf_1 rebuffer84 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ),
    .X(net116));
 sg13g2_buf_1 rebuffer85 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_mux2_1_A1_1_X ),
    .X(net117));
 sg13g2_buf_1 rebuffer86 (.A(net3182),
    .X(net118));
 sg13g2_buf_1 rebuffer87 (.A(\i_snitch.i_snitch_lsu.metadata_q[4]_sg13g2_o21ai_1_A1_B1_sg13g2_nand3_1_Y_B_sg13g2_and2_1_B_A_sg13g2_nand4_1_Y_D ),
    .X(net119));
 sg13g2_buf_1 rebuffer88 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_nand2_1_B_Y_sg13g2_and4_1_A_X ),
    .X(net120));
 sg13g2_buf_8 rebuffer89 (.A(net3181),
    .X(net121));
 sg13g2_buf_1 rebuffer90 (.A(net2536),
    .X(net122));
 sg13g2_buf_1 rebuffer91 (.A(net2608),
    .X(net123));
 sg13g2_buf_1 rebuffer92 (.A(net3128),
    .X(net124));
 sg13g2_buf_2 rebuffer93 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_full_q_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_B ),
    .X(net125));
 sg13g2_buf_1 rebuffer198 (.A(\i_snitch.pc_d[21]_sg13g2_a21oi_1_Y_B1_sg13g2_a221oi_1_Y_A2_sg13g2_xor2_1_X_B ),
    .X(net230));
 sg13g2_buf_16 rebuffer278 (.X(net310),
    .A(net2257));
 sg13g2_buf_1 rebuffer382 (.A(\i_snitch.pc_d[11]_sg13g2_a22oi_1_Y_B1_sg13g2_nand3_1_Y_C_sg13g2_or3_1_X_B_sg13g2_o21ai_1_A1_Y ),
    .X(net414));
 sg13g2_buf_1 rebuffer387 (.A(\i_snitch.pc_d[28]_sg13g2_a21oi_1_Y_B1 ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold391 (.A(data_pvalid),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[43]_sg13g2_dfrbpq_1_Q_D ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[45]_sg13g2_dfrbpq_1_Q_D ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[41]_sg13g2_dfrbpq_1_Q_D ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[44]_sg13g2_dfrbpq_1_Q_D ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[36]_sg13g2_dfrbpq_1_Q_D ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[34]_sg13g2_dfrbpq_1_Q_D ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[35]_sg13g2_dfrbpq_1_Q_D ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_snitch.i_snitch_regfile.mem[432] ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[37]_sg13g2_dfrbpq_1_Q_D ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp_sg13g2_a21o_1_X_B1_sg13g2_nor3_1_Y_A ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold410 (.A(\strb_reg_q[6] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold411 (.A(\strb_reg_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold412 (.A(\i_snitch.i_snitch_regfile.mem[225] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_snitch.i_snitch_regfile.mem[481] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold416 (.A(\cnt_q[2] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold417 (.A(\cnt_q[2]_sg13g2_a21oi_1_B1_Y ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold418 (.A(\cnt_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_snitch.i_snitch_regfile.mem[336] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_snitch.i_snitch_regfile.mem[193] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_snitch.i_snitch_regfile.mem[510] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_snitch.i_snitch_regfile.mem[446] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold423 (.A(\i_snitch.i_snitch_regfile.mem[430] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_snitch.i_snitch_regfile.mem[306] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_snitch.i_snitch_regfile.mem[353] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_snitch.i_snitch_regfile.mem[65] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold427 (.A(\strb_reg_q[3] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold428 (.A(\strb_reg_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold429 (.A(\shift_reg_q[15] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold430 (.A(\shift_reg_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold431 (.A(\i_snitch.i_snitch_regfile.mem[129] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_snitch.i_snitch_regfile.mem[161] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold433 (.A(\shift_reg_q[4] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold434 (.A(\shift_reg_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold435 (.A(\i_snitch.i_snitch_regfile.mem[377] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold436 (.A(\shift_reg_q[10] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold437 (.A(\shift_reg_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_snitch.i_snitch_regfile.mem[321] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold440 (.A(\strb_reg_q[4] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold441 (.A(\strb_reg_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold442 (.A(\shift_reg_q[5] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold443 (.A(\shift_reg_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold444 (.A(\shift_reg_q[13] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold445 (.A(\shift_reg_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_snitch.i_snitch_regfile.mem[112] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold447 (.A(\shift_reg_q[2] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold448 (.A(\shift_reg_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold449 (.A(\shift_reg_q[17] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold450 (.A(\shift_reg_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold451 (.A(\shift_reg_q[21] ),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold452 (.A(\shift_reg_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_snitch.i_snitch_regfile.mem[449] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold454 (.A(\shift_reg_q[14] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold455 (.A(\shift_reg_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_snitch.sb_q[4] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_snitch.sb_d[4]_sg13g2_o21ai_1_Y_B1 ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold458 (.A(\i_snitch.sb_q[15] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_snitch.sb_d[15]_sg13g2_o21ai_1_Y_B1 ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold460 (.A(\shift_reg_q[7] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold461 (.A(\shift_reg_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_snitch.i_snitch_regfile.mem[97] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_snitch.i_snitch_regfile.mem[385] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold464 (.A(\shift_reg_q[20] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold465 (.A(\shift_reg_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold466 (.A(\shift_reg_q[19] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold467 (.A(\shift_reg_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold468 (.A(\cnt_q[0] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold469 (.A(\strb_reg_q[0] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold470 (.A(\strb_reg_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold471 (.A(\shift_reg_q[8] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold472 (.A(\shift_reg_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_snitch.i_snitch_regfile.mem[257] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold474 (.A(\shift_reg_q[6] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold475 (.A(\shift_reg_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold476 (.A(\shift_reg_q[18] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold477 (.A(\shift_reg_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_snitch.i_snitch_regfile.mem[442] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold479 (.A(\shift_reg_q[23] ),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold480 (.A(\shift_reg_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_snitch.i_snitch_regfile.mem[458] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_snitch.i_snitch_regfile.mem[33] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold483 (.A(\shift_reg_q[25] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold484 (.A(\shift_reg_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold485 (.A(\strb_reg_q[2] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold486 (.A(\strb_reg_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold487 (.A(\shift_reg_q[11] ),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold488 (.A(\shift_reg_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold489 (.A(\shift_reg_q[3] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold490 (.A(\shift_reg_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_snitch.i_snitch_regfile.mem[80] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold492 (.A(\i_snitch.i_snitch_regfile.mem[417] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold493 (.A(\strb_reg_q[1] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold494 (.A(\strb_reg_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold495 (.A(\shift_reg_q[0] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold496 (.A(\shift_reg_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold497 (.A(\shift_reg_q[24] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold498 (.A(\shift_reg_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold499 (.A(\i_snitch.sb_q[8] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_snitch.sb_d[8]_sg13g2_o21ai_1_Y_B1 ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold502 (.A(\strb_reg_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_nor2_1_Y_A_sg13g2_and2_1_X_B ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold503 (.A(\shift_reg_q[1] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold504 (.A(\shift_reg_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold505 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold506 (.A(\shift_reg_q[9] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold507 (.A(\shift_reg_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_snitch.sb_q[5] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold509 (.A(\shift_reg_q[22] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold510 (.A(\shift_reg_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold511 (.A(\cnt_q[1] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_snitch.sb_q[7] ),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_snitch.wake_up_q[2] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold514 (.A(\shift_reg_q[16] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold515 (.A(\shift_reg_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold516 (.A(\shift_reg_q[12] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold517 (.A(\shift_reg_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold518 (.A(\shift_reg_q[26] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold519 (.A(\shift_reg_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold521 (.A(\i_snitch.wake_up_q[1] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_snitch.i_snitch_lsu.metadata_q[0] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_snitch.sb_q[12] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold524 (.A(\i_snitch.sb_d[12]_sg13g2_o21ai_1_Y_B1 ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_snitch.sb_q[13] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold526 (.A(\i_snitch.sb_d[13]_sg13g2_o21ai_1_Y_B1 ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold528 (.A(\i_snitch.sb_q[10] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_snitch.i_snitch_regfile.mem[273] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold531 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold532 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold533 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold534 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold535 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[38]_sg13g2_dfrbpq_1_Q_D ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold537 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_snitch.sb_q[9] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold539 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold541 (.A(\i_snitch.sb_q[11] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold542 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold544 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold546 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[39]_sg13g2_dfrbpq_1_Q_D ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold549 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold552 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold554 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold557 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold558 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold559 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold560 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold561 (.A(\i_snitch.sb_q[3] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold562 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold563 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_snitch.sb_q[6] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold565 (.A(\i_snitch.i_snitch_regfile.mem[415] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold567 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[32]_sg13g2_dfrbpq_1_Q_D ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_snitch.i_snitch_regfile.mem[325]_sg13g2_inv_1_A_Y ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold569 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold570 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold571 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold572 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold573 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold575 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold576 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[1] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold578 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold580 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold582 (.A(\shift_reg_q[27] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold583 (.A(\shift_reg_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold584 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold586 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[29] ),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold587 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold588 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold589 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold590 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[24] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold592 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[16]_sg13g2_dfrbpq_1_Q_D ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold594 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold596 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[40]_sg13g2_dfrbpq_1_Q_D ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[28] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold598 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold600 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9] ),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold602 (.A(\i_snitch.i_snitch_regfile.mem[264] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold604 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold606 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold607 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold608 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold609 (.A(\i_snitch.i_snitch_regfile.mem[324]_sg13g2_inv_1_A_Y ),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold610 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[4] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold611 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[0] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold612 (.A(\i_snitch.i_snitch_regfile.mem[265] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold614 (.A(\i_snitch.wake_up_q[0]_sg13g2_dfrbpq_1_Q_D_sg13g2_mux2_1_X_S_sg13g2_mux2_1_X_A1_sg13g2_nand2_1_Y_B_sg13g2_dfrbpq_1_Q_D ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold616 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold617 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold618 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold619 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold620 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold621 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold622 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold623 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[11] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold624 (.A(\i_snitch.i_snitch_regfile.mem[335] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold625 (.A(\i_snitch.i_snitch_regfile.mem[290]_sg13g2_inv_1_A_Y ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold626 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold627 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[33]_sg13g2_dfrbpq_1_Q_D ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold628 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold629 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[42]_sg13g2_dfrbpq_1_Q_D ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold630 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold631 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold632 (.A(\i_snitch.i_snitch_regfile.mem[328] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold633 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[5] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold634 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold635 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[14] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold636 (.A(\i_snitch.sb_q[2] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold637 (.A(\i_snitch.inst_addr_o[1] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold638 (.A(\i_snitch.i_snitch_regfile.mem[283] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold639 (.A(\i_snitch.i_snitch_regfile.mem[286] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_snitch.i_snitch_regfile.mem[338] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold641 (.A(\i_snitch.i_snitch_regfile.mem[261]_sg13g2_inv_1_A_Y ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold642 (.A(\i_snitch.i_snitch_regfile.mem[389]_sg13g2_inv_1_A_Y ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold643 (.A(\i_snitch.i_snitch_regfile.mem[451]_sg13g2_inv_1_A_Y ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold644 (.A(\data_pdata[5] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold645 (.A(\data_pdata[5]_sg13g2_dfrbpq_1_Q_D ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_snitch.i_snitch_regfile.mem[291]_sg13g2_inv_1_A_Y ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold647 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold648 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.b_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold649 (.A(\data_pdata[7] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold650 (.A(\data_pdata[7]_sg13g2_dfrbpq_1_Q_D ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold651 (.A(\i_snitch.i_snitch_regfile.mem[282] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold652 (.A(\data_pdata[0] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold653 (.A(\data_pdata[0]_sg13g2_dfrbpq_1_Q_D ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold654 (.A(\data_pdata[2] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold655 (.A(\data_pdata[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold656 (.A(\data_pdata[3] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold657 (.A(\data_pdata[3]_sg13g2_dfrbpq_1_Q_D ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold658 (.A(\i_snitch.i_snitch_regfile.mem[322]_sg13g2_inv_1_A_Y ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold659 (.A(\i_snitch.i_snitch_regfile.mem[277] ),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold660 (.A(\i_snitch.i_snitch_lsu.metadata_q[9] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_snitch.i_snitch_regfile.mem[260]_sg13g2_inv_1_A_Y ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold662 (.A(\i_snitch.i_snitch_regfile.mem[387]_sg13g2_inv_1_A_Y ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold663 (.A(\i_snitch.sb_q[1] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold664 (.A(\i_snitch.inst_addr_o[31] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold665 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[27] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold666 (.A(\data_pdata[4] ),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold667 (.A(\data_pdata[4]_sg13g2_dfrbpq_1_Q_D ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold668 (.A(\i_snitch.i_snitch_regfile.mem[281] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold669 (.A(\i_snitch.i_snitch_regfile.mem[258]_sg13g2_inv_1_A_Y ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold670 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[21] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold671 (.A(\i_snitch.i_snitch_regfile.mem[346] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_snitch.i_snitch_regfile.mem[269] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold673 (.A(\i_snitch.i_snitch_regfile.mem[172] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold674 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15]_sg13g2_dfrbpq_1_Q_D ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold676 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[12] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold677 (.A(\i_snitch.i_snitch_regfile.mem[331] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold678 (.A(\i_snitch.sb_q[14] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold679 (.A(\i_snitch.sb_d[14]_sg13g2_o21ai_1_Y_B1 ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold680 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold681 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24]_sg13g2_dfrbpq_1_Q_D ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold682 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[31] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold683 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[23] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold684 (.A(\i_snitch.i_snitch_regfile.mem[471] ),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_snitch.i_snitch_regfile.mem[320] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold686 (.A(\i_snitch.i_snitch_regfile.mem[212] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold687 (.A(\data_pdata[6] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold688 (.A(\data_pdata[6]_sg13g2_dfrbpq_1_Q_D ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold689 (.A(\data_pdata[23] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold690 (.A(\data_pdata[23]_sg13g2_dfrbpq_1_Q_D ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold691 (.A(\i_snitch.i_snitch_regfile.mem[337] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold692 (.A(\i_snitch.i_snitch_regfile.mem[244] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold693 (.A(\data_pdata[13] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold694 (.A(\data_pdata[13]_sg13g2_dfrbpq_1_Q_D ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold695 (.A(\i_snitch.i_snitch_regfile.mem[177] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold696 (.A(\i_snitch.i_snitch_regfile.mem[127] ),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold697 (.A(\data_pdata[17] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold698 (.A(\data_pdata[17]_sg13g2_dfrbpq_1_Q_D ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold699 (.A(\i_snitch.i_snitch_regfile.mem[95] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold700 (.A(\i_snitch.i_snitch_regfile.mem[152] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold701 (.A(\i_snitch.i_snitch_regfile.mem[329] ),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold702 (.A(\data_pdata[1] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold703 (.A(\data_pdata[1]_sg13g2_dfrbpq_1_Q_D ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold704 (.A(\i_snitch.i_snitch_regfile.mem[105] ),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold705 (.A(\i_snitch.i_snitch_regfile.mem[360] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold706 (.A(\i_snitch.i_snitch_regfile.mem[137] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold707 (.A(\i_snitch.i_snitch_regfile.mem[201] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold708 (.A(\i_snitch.i_snitch_regfile.mem[140] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_snitch.i_snitch_regfile.mem[128] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold710 (.A(\i_snitch.i_snitch_regfile.mem[448] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold711 (.A(\i_snitch.i_snitch_regfile.mem[342] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold712 (.A(\i_snitch.i_snitch_regfile.mem[463] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold713 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold714 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19]_sg13g2_dfrbpq_1_Q_D ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold715 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0] ),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold716 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[0]_sg13g2_dfrbpq_1_Q_D ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold717 (.A(\data_pdata[18] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold718 (.A(\data_pdata[18]_sg13g2_dfrbpq_1_Q_D ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold719 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[2] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold720 (.A(\i_snitch.i_snitch_regfile.mem[136] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold721 (.A(\i_snitch.i_snitch_regfile.mem[374] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold722 (.A(\data_pdata[19] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold723 (.A(\data_pdata[19]_sg13g2_dfrbpq_1_Q_D ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold724 (.A(\i_snitch.i_snitch_regfile.mem[223] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold725 (.A(\i_snitch.i_snitch_regfile.mem[439] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold726 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26]_sg13g2_dfrbpq_1_Q_D ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold728 (.A(\i_snitch.i_snitch_regfile.mem[392] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold729 (.A(\i_snitch.i_snitch_regfile.mem[255] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold730 (.A(\i_snitch.i_snitch_regfile.mem[460] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold731 (.A(\i_req_arb.gen_arbiter.rr_q ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold732 (.A(\i_req_arb.gen_arbiter.rr_q_sg13g2_a22oi_1_A1_Y ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold733 (.A(\i_snitch.i_snitch_regfile.mem[64] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold734 (.A(\i_snitch.i_snitch_regfile.mem[88] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold735 (.A(\i_snitch.i_snitch_regfile.mem[145] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold736 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[45] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold737 (.A(\i_snitch.i_snitch_regfile.mem[86] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold738 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold739 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8]_sg13g2_dfrbpq_1_Q_D ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold740 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold741 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7]_sg13g2_dfrbpq_1_Q_D ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold742 (.A(\i_snitch.i_snitch_regfile.mem[465] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold743 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold744 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30]_sg13g2_dfrbpq_1_Q_D ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold745 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold746 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29]_sg13g2_dfrbpq_1_Q_D ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold747 (.A(\i_snitch.i_snitch_regfile.mem[425] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold748 (.A(\i_snitch.i_snitch_regfile.mem[388]_sg13g2_inv_1_A_Y ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold749 (.A(\i_snitch.i_snitch_regfile.mem[345] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold750 (.A(\i_snitch.i_snitch_regfile.mem[251] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_snitch.i_snitch_regfile.mem[224] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold752 (.A(\i_snitch.i_snitch_regfile.mem[503] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold753 (.A(\i_snitch.i_snitch_regfile.mem[276] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold754 (.A(\i_snitch.i_snitch_regfile.mem[326] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold755 (.A(\i_snitch.i_snitch_regfile.mem[267] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold756 (.A(\i_snitch.i_snitch_regfile.mem[457] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold757 (.A(\i_snitch.i_snitch_regfile.mem[479] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold758 (.A(\i_snitch.i_snitch_regfile.mem[184] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold759 (.A(\i_snitch.i_snitch_regfile.mem[215] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold760 (.A(\i_snitch.i_snitch_regfile.mem[433] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold761 (.A(\i_snitch.i_snitch_regfile.mem[399] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold762 (.A(\i_snitch.i_snitch_regfile.mem[73] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold763 (.A(\i_snitch.i_snitch_regfile.mem[361] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold764 (.A(\i_snitch.i_snitch_regfile.mem[440] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold765 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[20] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold766 (.A(\data_pdata[22] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold767 (.A(\data_pdata[22]_sg13g2_dfrbpq_1_Q_D ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold768 (.A(\i_snitch.i_snitch_regfile.mem[393] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold769 (.A(\i_snitch.i_snitch_regfile.mem[438] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold770 (.A(\i_snitch.i_snitch_regfile.mem[383] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold771 (.A(\data_pdata[21] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold772 (.A(\data_pdata[21]_sg13g2_dfrbpq_1_Q_D ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold773 (.A(\i_snitch.i_snitch_regfile.mem[429] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold774 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28]_sg13g2_dfrbpq_1_Q_D ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold776 (.A(\i_snitch.i_snitch_regfile.mem[216] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold777 (.A(\data_pdata[16] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold778 (.A(\data_pdata[16]_sg13g2_dfrbpq_1_Q_D ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_snitch.i_snitch_regfile.mem[268] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold780 (.A(\i_snitch.i_snitch_regfile.mem[63] ),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold781 (.A(\i_snitch.i_snitch_regfile.mem[351] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_snitch.i_snitch_regfile.mem[76] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold783 (.A(\i_snitch.i_snitch_regfile.mem[456] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold784 (.A(\i_snitch.i_snitch_regfile.mem[424] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold785 (.A(\i_snitch.i_snitch_regfile.mem[107] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold786 (.A(\data_pdata[26] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold787 (.A(\data_pdata[26]_sg13g2_dfrbpq_1_Q_D ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold788 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold789 (.A(\i_snitch.i_snitch_regfile.mem[40] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold790 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[13] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold791 (.A(\i_snitch.i_snitch_regfile.mem[200] ),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold792 (.A(\data_pdata[10] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold793 (.A(\data_pdata[10]_sg13g2_dfrbpq_1_Q_D ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold794 (.A(\i_snitch.i_snitch_regfile.mem[475] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold795 (.A(\i_snitch.i_snitch_regfile.mem[408] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold796 (.A(\i_snitch.i_snitch_regfile.mem[146] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold797 (.A(\i_snitch.i_snitch_regfile.mem[431] ),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold798 (.A(\i_snitch.i_snitch_regfile.mem[57] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold799 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold800 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31]_sg13g2_dfrbpq_1_Q_D ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold801 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold802 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21]_sg13g2_dfrbpq_1_Q_D ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold803 (.A(\i_snitch.i_snitch_regfile.mem[238] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold804 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold805 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23]_sg13g2_dfrbpq_1_Q_D ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_snitch.i_snitch_regfile.mem[473] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold807 (.A(\i_snitch.i_snitch_regfile.mem[364] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold808 (.A(\i_snitch.i_snitch_regfile.mem[191] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold809 (.A(\i_snitch.i_snitch_regfile.mem[41] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold810 (.A(\i_snitch.i_snitch_regfile.mem[511] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold811 (.A(\i_snitch.i_snitch_regfile.mem[111] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold812 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[43] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold813 (.A(\i_snitch.i_snitch_regfile.mem[47] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold814 (.A(\data_pdata[29] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold815 (.A(\data_pdata[29]_sg13g2_dfrbpq_1_Q_D ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold816 (.A(\i_snitch.i_snitch_regfile.mem[363] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold817 (.A(\i_snitch.i_snitch_regfile.mem[104] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold818 (.A(\i_snitch.i_snitch_regfile.mem[397] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold819 (.A(\i_snitch.i_snitch_regfile.mem[151] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold820 (.A(\i_snitch.i_snitch_regfile.mem[138] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold821 (.A(\i_snitch.i_snitch_regfile.mem[150] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold822 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold823 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18]_sg13g2_dfrbpq_1_Q_D ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold824 (.A(\i_snitch.i_snitch_regfile.mem[454] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_snitch.i_snitch_regfile.mem[217] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold826 (.A(\data_pdata[31] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold827 (.A(\data_pdata[31]_sg13g2_dfrbpq_1_Q_D ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold828 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[44] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_snitch.i_snitch_regfile.mem[32] ),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold830 (.A(\i_snitch.i_snitch_regfile.mem[472] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold831 (.A(\i_snitch.i_snitch_regfile.mem[211] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold832 (.A(\i_snitch.i_snitch_regfile.mem[340] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold833 (.A(\i_snitch.i_snitch_regfile.mem[256] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold834 (.A(\i_snitch.i_snitch_regfile.mem[180] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold835 (.A(\i_snitch.i_snitch_regfile.mem[53] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold836 (.A(\i_snitch.i_snitch_regfile.mem[504] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold837 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[6] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold838 (.A(\i_snitch.i_snitch_regfile.mem[203] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold839 (.A(\i_snitch.i_snitch_regfile.mem[148] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold840 (.A(\i_snitch.i_snitch_regfile.mem[96] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold841 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold842 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11]_sg13g2_dfrbpq_1_Q_D ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold843 (.A(\i_snitch.i_snitch_regfile.mem[489] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold844 (.A(\i_snitch.i_snitch_regfile.mem[94] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold845 (.A(\i_snitch.i_snitch_regfile.mem[85] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold846 (.A(\i_snitch.i_snitch_regfile.mem[486] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold847 (.A(\i_snitch.i_snitch_regfile.mem[344] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold848 (.A(\i_snitch.i_snitch_regfile.mem[52] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold849 (.A(\i_snitch.i_snitch_regfile.mem[470] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold850 (.A(\i_snitch.i_snitch_regfile.mem[488] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold851 (.A(\i_snitch.i_snitch_regfile.mem[395] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold852 (.A(\i_snitch.i_snitch_regfile.mem[285] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold853 (.A(\i_snitch.i_snitch_regfile.mem[199] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold854 (.A(\i_snitch.i_snitch_regfile.mem[416] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_snitch.i_snitch_regfile.mem[155] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold856 (.A(\i_snitch.i_snitch_regfile.mem[369] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold857 (.A(\data_pdata[9] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold858 (.A(\data_pdata[9]_sg13g2_dfrbpq_1_Q_D ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_snitch.i_snitch_regfile.mem[343] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold860 (.A(\i_snitch.i_snitch_regfile.mem[459] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold861 (.A(\i_snitch.inst_addr_o[17] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold862 (.A(\i_snitch.i_snitch_regfile.mem[347] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold863 (.A(\i_snitch.i_snitch_regfile.mem[367] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold864 (.A(\i_snitch.i_snitch_regfile.mem[235] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold865 (.A(\i_snitch.i_snitch_regfile.mem[171] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_snitch.i_snitch_regfile.mem[407] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold867 (.A(\i_snitch.i_snitch_regfile.mem[248] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold868 (.A(\i_snitch.i_snitch_regfile.mem[72] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold869 (.A(\data_pdata[12] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold870 (.A(\data_pdata[12]_sg13g2_dfrbpq_1_Q_D ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold871 (.A(\i_snitch.i_snitch_regfile.mem[246] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold872 (.A(\i_snitch.i_snitch_regfile.mem[375] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold873 (.A(\i_snitch.i_snitch_regfile.mem[468] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold874 (.A(\i_snitch.i_snitch_regfile.mem[175] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold875 (.A(\rsp_data_q[20] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold876 (.A(\rsp_data_q[20]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold877 (.A(\i_snitch.i_snitch_regfile.mem[348] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold878 (.A(\i_snitch.i_snitch_regfile.mem[160] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold879 (.A(\i_snitch.i_snitch_regfile.mem[110] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold880 (.A(\i_snitch.i_snitch_regfile.mem[279] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold881 (.A(\i_snitch.i_snitch_regfile.mem[202] ),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold882 (.A(rsp_state_q),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold883 (.A(target_sel_q_sg13g2_nand2b_1_A_N_Y),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q_sg13g2_dfrbpq_1_Q_D ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold885 (.A(\i_snitch.i_snitch_regfile.mem[287] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold886 (.A(\i_snitch.i_snitch_regfile.mem[230] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold887 (.A(\i_snitch.i_snitch_regfile.mem[74] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold888 (.A(\i_snitch.i_snitch_regfile.mem[56] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold889 (.A(\i_snitch.i_snitch_regfile.mem[254] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold890 (.A(\i_snitch.i_snitch_regfile.mem[113] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold891 (.A(\i_snitch.i_snitch_regfile.mem[61] ),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold892 (.A(\i_snitch.i_snitch_regfile.mem[159] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold893 (.A(\data_pdata[20] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold894 (.A(\i_snitch.i_snitch_regfile.mem[204] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold895 (.A(\data_pdata[24] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold896 (.A(\data_pdata[24]_sg13g2_dfrbpq_1_Q_D ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold897 (.A(\i_snitch.i_snitch_regfile.mem[83] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold898 (.A(\i_snitch.i_snitch_regfile.mem[362] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold899 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[41] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold900 (.A(\i_snitch.i_snitch_regfile.mem[477] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold901 (.A(\i_snitch.i_snitch_regfile.mem[447] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold902 (.A(\i_snitch.i_snitch_regfile.mem[75] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold903 (.A(\i_snitch.i_snitch_regfile.mem[478] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold904 (.A(\i_snitch.i_snitch_regfile.mem[428] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold905 (.A(\i_snitch.i_snitch_regfile.mem[156] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold906 (.A(\i_snitch.i_snitch_regfile.mem[135] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold907 (.A(\i_snitch.i_snitch_regfile.mem[87] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold908 (.A(\i_snitch.i_snitch_regfile.mem[270] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold909 (.A(\data_pdata[27] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold910 (.A(\data_pdata[27]_sg13g2_dfrbpq_1_Q_D ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold911 (.A(\i_snitch.i_snitch_regfile.mem[469] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold912 (.A(\i_snitch.i_snitch_regfile.mem[278] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold913 (.A(\data_pdata[25] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold914 (.A(\data_pdata[25]_sg13g2_dfrbpq_1_Q_D ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold915 (.A(\i_snitch.i_snitch_regfile.mem[334] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold916 (.A(\i_snitch.i_snitch_regfile.mem[341] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold917 (.A(\i_snitch.i_snitch_regfile.mem[332] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold918 (.A(\rsp_data_q[16] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold919 (.A(\rsp_data_q[16]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold920 (.A(\i_snitch.i_snitch_regfile.mem[494] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold921 (.A(\i_snitch.i_snitch_regfile.mem[168] ),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold922 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold923 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[1]_sg13g2_dfrbpq_1_Q_D ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold924 (.A(\i_snitch.i_snitch_regfile.mem[497] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold925 (.A(\i_snitch.i_snitch_regfile.mem[352] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold926 (.A(\i_snitch.i_snitch_regfile.mem[253] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_snitch.i_snitch_regfile.mem[141] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold928 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold929 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[2]_sg13g2_dfrbpq_1_Q_D ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold930 (.A(\i_snitch.i_snitch_regfile.mem[89] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold931 (.A(\i_snitch.i_snitch_regfile.mem[327] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold932 (.A(\i_snitch.i_snitch_regfile.mem[350] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold933 (.A(\i_snitch.i_snitch_regfile.mem[134] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold934 (.A(\data_pdata[15] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold935 (.A(\data_pdata[15]_sg13g2_dfrbpq_1_Q_D ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold936 (.A(\i_snitch.i_snitch_regfile.mem[210] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold937 (.A(\i_snitch.i_snitch_regfile.mem[500] ),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold938 (.A(\i_snitch.i_snitch_regfile.mem[220] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold939 (.A(\i_snitch.i_snitch_regfile.mem[158] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold940 (.A(\i_snitch.i_snitch_regfile.mem[222] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold941 (.A(\i_snitch.i_snitch_regfile.mem[480] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold942 (.A(\i_snitch.i_snitch_regfile.mem[174] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold943 (.A(\i_snitch.i_snitch_regfile.mem[401] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold944 (.A(\i_snitch.i_snitch_regfile.mem[333] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold945 (.A(\i_snitch.i_snitch_regfile.mem[79] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold946 (.A(\i_snitch.i_snitch_regfile.mem[51] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold947 (.A(\i_snitch.i_snitch_regfile.mem[241] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold948 (.A(\i_snitch.i_snitch_regfile.mem[208] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold949 (.A(\i_snitch.i_snitch_regfile.mem[58] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold950 (.A(\i_snitch.i_snitch_regfile.mem[118] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold951 (.A(\i_snitch.i_snitch_regfile.mem[464] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold952 (.A(\i_snitch.i_snitch_regfile.mem[219] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold953 (.A(\i_snitch.i_snitch_regfile.mem[372] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold954 (.A(\i_snitch.i_snitch_regfile.mem[370] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold955 (.A(\i_snitch.i_snitch_regfile.mem[71] ),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold956 (.A(\i_snitch.i_snitch_regfile.mem[371] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold957 (.A(\i_snitch.i_snitch_regfile.mem[274] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold958 (.A(\i_snitch.inst_addr_o[10] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold959 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold960 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9]_sg13g2_dfrbpq_1_Q_D ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold961 (.A(\i_snitch.i_snitch_regfile.mem[250] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold962 (.A(\i_snitch.i_snitch_regfile.mem[84] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold963 (.A(\data_pdata[11] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold964 (.A(\data_pdata[11]_sg13g2_dfrbpq_1_Q_D ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold965 (.A(\i_snitch.i_snitch_regfile.mem[330] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold966 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold967 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5]_sg13g2_dfrbpq_1_Q_D ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold968 (.A(\i_snitch.i_snitch_regfile.mem[379] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold969 (.A(\i_snitch.i_snitch_regfile.mem[495] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold970 (.A(\i_snitch.i_snitch_regfile.mem[173] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold971 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold972 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold973 (.A(\i_snitch.i_snitch_regfile.mem[247] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold974 (.A(\i_snitch.i_snitch_regfile.mem[249] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold975 (.A(\i_snitch.i_snitch_regfile.mem[109] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold976 (.A(\i_snitch.i_snitch_regfile.mem[455] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold977 (.A(\i_snitch.i_snitch_regfile.mem[154] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold978 (.A(\i_snitch.i_snitch_regfile.mem[82] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold979 (.A(\i_snitch.i_snitch_regfile.mem[60] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold980 (.A(\i_snitch.i_snitch_regfile.mem[242] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold981 (.A(\i_snitch.i_snitch_regfile.mem[38] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold982 (.A(\i_snitch.i_snitch_regfile.mem[365] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold983 (.A(\i_snitch.i_snitch_regfile.mem[108] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold984 (.A(\i_snitch.i_snitch_regfile.mem[221] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold985 (.A(\i_snitch.i_snitch_regfile.mem[493] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold986 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold987 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[4]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold988 (.A(\i_snitch.i_snitch_regfile.mem[266] ),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold989 (.A(\i_snitch.i_snitch_regfile.mem[378] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold990 (.A(\i_snitch.i_snitch_regfile.mem[381] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold991 (.A(\i_snitch.i_snitch_regfile.mem[243] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i_snitch.i_snitch_regfile.mem[252] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold993 (.A(\i_snitch.i_snitch_regfile.mem[491] ),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold994 (.A(target_sel_q),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold995 (.A(target_sel_q_sg13g2_dfrbpq_1_Q_D),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold996 (.A(\i_snitch.i_snitch_regfile.mem[234] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold997 (.A(\i_snitch.i_snitch_regfile.mem[169] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold998 (.A(\i_snitch.i_snitch_regfile.mem[271] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold999 (.A(\i_snitch.i_snitch_regfile.mem[359] ),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\i_snitch.i_snitch_regfile.mem[233] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\i_snitch.i_snitch_regfile.mem[147] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\i_snitch.i_snitch_regfile.mem[436] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\data_pdata[14] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\data_pdata[14]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\i_snitch.i_snitch_regfile.mem[92] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\i_snitch.i_snitch_regfile.mem[91] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold1007 (.A(\i_snitch.i_snitch_regfile.mem[209] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\i_snitch.i_snitch_regfile.mem[62] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\i_snitch.i_snitch_regfile.mem[205] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\i_snitch.i_snitch_regfile.mem[461] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\i_snitch.i_snitch_regfile.mem[182] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\i_snitch.i_snitch_regfile.mem[45] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\i_snitch.i_snitch_regfile.mem[144] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\i_snitch.i_snitch_regfile.mem[192] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold1018 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\rsp_data_q[28] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\rsp_data_q[28]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\i_snitch.i_snitch_regfile.mem[39] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\data_pdata[30] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\data_pdata[30]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\i_snitch.i_snitch_regfile.mem[236] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\i_snitch.i_snitch_regfile.mem[49] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\i_snitch.i_snitch_regfile.mem[240] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\i_snitch.i_snitch_regfile.mem[119] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\i_snitch.i_snitch_regfile.mem[116] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[22] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\i_snitch.i_snitch_regfile.mem[231] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\i_snitch.i_snitch_regfile.mem[284] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\i_snitch.i_snitch_regfile.mem[427] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\i_snitch.i_snitch_regfile.mem[339] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\i_snitch.i_snitch_regfile.mem[59] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\i_snitch.i_snitch_regfile.mem[102] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\i_snitch.i_snitch_regfile.mem[349] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\i_req_arb.data_i[44] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\i_snitch.inst_addr_o[27] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\i_snitch.i_snitch_regfile.mem[50] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\i_snitch.i_snitch_regfile.mem[384] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\i_snitch.i_snitch_regfile.mem[183] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_snitch.i_snitch_regfile.mem[43] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold1048 (.A(\i_snitch.i_snitch_regfile.mem[207] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\i_snitch.i_snitch_regfile.mem[303] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\i_snitch.i_snitch_regfile.mem[44] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\data_pdata[28] ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold1052 (.A(\i_snitch.i_snitch_regfile.mem[206] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\i_snitch.i_snitch_regfile.mem[149] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\i_snitch.i_snitch_regfile.mem[120] ),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\i_snitch.i_snitch_regfile.mem[78] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\i_snitch.i_snitch_regfile.mem[218] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.b_data_q[3] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\i_snitch.i_snitch_regfile.mem[368] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\i_snitch.i_snitch_regfile.mem[245] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\i_snitch.i_snitch_regfile.mem[462] ),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\i_snitch.i_snitch_regfile.mem[139] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\i_snitch.i_snitch_regfile.mem[157] ),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\i_snitch.i_snitch_regfile.mem[474] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\i_snitch.i_snitch_regfile.mem[406] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\i_snitch.i_snitch_regfile.mem[422] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\i_snitch.i_snitch_regfile.mem[358] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\i_snitch.i_snitch_regfile.mem[70] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold1074 (.A(\i_snitch.i_snitch_regfile.mem[214] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\rsp_data_q[31] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\rsp_data_q[31]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\i_snitch.i_snitch_regfile.mem[502] ),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\i_snitch.i_snitch_regfile.mem[90] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\i_snitch.i_snitch_regfile.mem[404] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\i_snitch.i_snitch_regfile.mem[492] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\i_snitch.i_snitch_regfile.mem[198] ),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\i_snitch.i_snitch_regfile.mem[263] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\i_snitch.i_snitch_regfile.mem[77] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\i_snitch.i_snitch_regfile.mem[142] ),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\i_snitch.i_snitch_regfile.mem[54] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\i_snitch.i_snitch_regfile.mem[280] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\i_req_arb.data_i[38] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_snitch.i_snitch_regfile.mem[476] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\i_snitch.i_snitch_regfile.mem[396] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\i_snitch.wake_up_q[0] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\i_snitch.i_snitch_regfile.mem[466] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\i_snitch.i_snitch_regfile.mem[46] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\i_snitch.i_snitch_regfile.mem[382] ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\i_snitch.i_snitch_regfile.mem[239] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\i_snitch.i_snitch_regfile.mem[412] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\i_snitch.i_snitch_regfile.mem[398] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\i_snitch.i_snitch_regfile.mem[93] ),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\i_snitch.i_snitch_regfile.mem[213] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\i_snitch.i_snitch_regfile.mem[166] ),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\i_snitch.i_snitch_regfile.mem[506] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\i_snitch.i_snitch_regfile.mem[232] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\i_snitch.i_snitch_regfile.mem[300] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3] ),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[3]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\i_snitch.i_snitch_regfile.mem[373] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\i_snitch.i_snitch_regfile.mem[143] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\i_snitch.i_snitch_regfile.mem[275] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\i_snitch.i_snitch_regfile.mem[237] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_snitch.i_snitch_regfile.mem[390] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\i_snitch.i_snitch_regfile.mem[434] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\data_pdata[8] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\data_pdata[8]_sg13g2_dfrbpq_1_Q_D ),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[39] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\i_snitch.i_snitch_regfile.mem[262] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\i_snitch.i_snitch_regfile.mem[153] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\i_snitch.i_snitch_regfile.mem[310] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\rsp_data_q[15] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\rsp_data_q[15]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\i_snitch.i_snitch_regfile.mem[414] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[14] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\rsp_data_q[30] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\rsp_data_q[30]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\i_snitch.i_snitch_regfile.mem[467] ),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\i_snitch.i_snitch_lsu.metadata_q[4] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\i_snitch.i_snitch_regfile.mem[318] ),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\i_snitch.i_snitch_regfile.mem[315] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\i_snitch.i_snitch_regfile.mem[167] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\i_snitch.i_snitch_regfile.mem[402] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\i_snitch.i_snitch_regfile.mem[115] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\i_snitch.inst_addr_o[19] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\rsp_data_q[24] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\i_snitch.i_snitch_regfile.mem[42] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\rsp_data_q[22] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\rsp_data_q[22]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\i_snitch.i_snitch_regfile.mem[316] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_snitch.i_snitch_regfile.mem[121] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold1141 (.A(\i_snitch.i_snitch_regfile.mem[380] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\i_snitch.consec_pc[0] ),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\i_snitch.i_snitch_regfile.mem[181] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\i_snitch.i_snitch_regfile.mem[411] ),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[12] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\i_snitch.i_snitch_regfile.mem[178] ),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\i_snitch.i_snitch_regfile.mem[409] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\i_snitch.i_snitch_regfile.mem[125] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[36] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\i_snitch.i_snitch_regfile.mem[311] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\rsp_data_q[8] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\rsp_data_q[8]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\i_snitch.i_snitch_regfile.mem[426] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_snitch.i_snitch_regfile.mem[441] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\i_snitch.i_snitch_regfile.mem[185] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\i_snitch.i_snitch_regfile.mem[501] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\i_snitch.i_snitch_regfile.mem[188] ),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\i_snitch.i_snitch_regfile.mem[376] ),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\i_snitch.i_snitch_regfile.mem[170] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[10] ),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\i_snitch.i_snitch_regfile.mem[366] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_snitch.i_snitch_regfile.mem[308] ),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold1164 (.A(\i_req_arb.data_i[42] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_snitch.inst_addr_o[25] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\i_snitch.i_snitch_regfile.mem[48] ),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\i_snitch.i_snitch_regfile.mem[505] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[17] ),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\i_snitch.i_snitch_regfile.mem[124] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\i_snitch.i_snitch_regfile.mem[444] ),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\i_snitch.i_snitch_regfile.mem[81] ),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\i_snitch.i_snitch_regfile.mem[117] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_snitch.i_snitch_regfile.mem[314] ),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold1174 (.A(\i_snitch.i_snitch_regfile.mem[355] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[25] ),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[8] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\i_snitch.i_snitch_regfile.mem[294] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[7] ),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\i_snitch.i_snitch_regfile.mem[317] ),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[31] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[9] ),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\i_snitch.i_snitch_regfile.mem[445] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\i_snitch.i_snitch_regfile.mem[186] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\i_snitch.i_snitch_regfile.mem[126] ),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[32] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\i_snitch.i_snitch_regfile.mem[295] ),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\i_snitch.i_snitch_regfile.mem[67] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\i_snitch.i_snitch_regfile.mem[405] ),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\i_snitch.i_snitch_regfile.mem[309] ),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\i_snitch.i_snitch_regfile.mem[507] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\rsp_data_q[11] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\rsp_data_q[11]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\i_snitch.i_snitch_regfile.mem[400] ),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\rsp_data_q[18] ),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\rsp_data_q[18]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[26] ),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\i_snitch.i_snitch_regfile.mem[272] ),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[29] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\i_snitch.i_snitch_regfile.mem[302] ),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\i_snitch.i_snitch_regfile.mem[319] ),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[24] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\i_snitch.i_snitch_regfile.mem[123] ),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\i_req_arb.data_i[40] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[42] ),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_snitch.i_snitch_regfile.mem[68] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold1206 (.A(\i_snitch.i_snitch_regfile.mem[194] ),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\i_snitch.i_snitch_regfile.mem[165] ),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[18] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\i_snitch.i_snitch_regfile.mem[490] ),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\i_snitch.inst_addr_o[21] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_snitch.i_snitch_regfile.mem[304] ),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\i_snitch.i_snitch_regfile.mem[190] ),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\i_snitch.gpr_waddr[4] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\i_snitch.i_snitch_regfile.mem[312] ),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\i_snitch.i_snitch_regfile.mem[132] ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\i_snitch.i_snitch_regfile.mem[496] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\i_snitch.i_snitch_regfile.mem[485] ),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\i_snitch.i_snitch_regfile.mem[122] ),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\i_snitch.i_snitch_regfile.mem[394] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[34] ),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[40] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\i_snitch.i_snitch_regfile.mem[288] ),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\i_snitch.i_snitch_regfile.mem[435] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\i_snitch.i_snitch_lsu.metadata_q[1] ),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\i_snitch.i_snitch_regfile.mem[298] ),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[11] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_snitch.i_snitch_regfile.mem[179] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\i_snitch.i_snitch_regfile.mem[301] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\i_snitch.i_snitch_regfile.mem[498] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\i_snitch.i_snitch_regfile.mem[410] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\rsp_data_q[4] ),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\rsp_data_q[4]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[33] ),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\i_snitch.i_snitch_regfile.mem[305] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\i_snitch.i_snitch_regfile.mem[509] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\i_snitch.i_snitch_regfile.mem[313] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[37] ),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\i_snitch.i_snitch_regfile.mem[450] ),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\rsp_data_q[23] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\rsp_data_q[23]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\i_snitch.i_snitch_regfile.mem[114] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[28] ),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\i_snitch.i_snitch_regfile.mem[176] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\i_snitch.i_snitch_regfile.mem[189] ),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\i_snitch.i_snitch_regfile.mem[483] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\i_snitch.i_snitch_regfile.mem[187] ),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\i_snitch.i_snitch_regfile.mem[35] ),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\i_snitch.i_snitch_regfile.mem[297] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\i_snitch.i_snitch_regfile.mem[452] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\i_snitch.i_snitch_regfile.mem[162] ),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[19] ),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\i_snitch.i_snitch_regfile.mem[356] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\i_snitch.i_snitch_regfile.mem[443] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\i_snitch.i_snitch_regfile.mem[130] ),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold1255 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[16] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\i_snitch.i_snitch_regfile.mem[69] ),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\i_snitch.i_snitch_regfile.mem[131] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\i_snitch.i_snitch_regfile.mem[164] ),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[21] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\i_snitch.i_snitch_regfile.mem[307] ),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\rsp_data_q[29] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\rsp_data_q[29]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_snitch.i_snitch_regfile.mem[103] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\i_snitch.i_snitch_regfile.mem[437] ),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\rsp_data_q[14] ),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\rsp_data_q[14]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\rsp_data_q[7] ),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\rsp_data_q[7]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\i_snitch.i_snitch_regfile.mem[419] ),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\i_snitch.i_snitch_regfile.mem[106] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[22] ),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\i_snitch.i_snitch_regfile.mem[293] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\i_snitch.i_snitch_regfile.mem[100] ),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\rsp_data_q[12] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\i_snitch.i_snitch_regfile.mem[482] ),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\i_snitch.i_snitch_regfile.mem[413] ),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\i_snitch.i_snitch_regfile.mem[163] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[13] ),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\i_snitch.i_snitch_regfile.mem[323] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\i_snitch.i_snitch_regfile.mem[197] ),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\i_snitch.i_snitch_regfile.mem[484] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\i_snitch.i_snitch_regfile.mem[487] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\i_snitch.i_snitch_regfile.mem[420] ),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\i_snitch.i_snitch_regfile.mem[289] ),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\i_snitch.i_snitch_regfile.mem[391] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\i_snitch.i_snitch_regfile.mem[296] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\i_snitch.i_snitch_regfile.mem[292] ),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\i_snitch.i_snitch_regfile.mem[453] ),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\rsp_data_q[6] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\rsp_data_q[6]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\i_snitch.i_snitch_regfile.mem[508] ),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\i_snitch.i_snitch_regfile.mem[499] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\i_snitch.i_snitch_regfile.mem[34] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\i_snitch.i_snitch_regfile.mem[227] ),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\i_snitch.i_snitch_regfile.mem[421] ),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\i_snitch.i_snitch_regfile.mem[196] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\rsp_data_q[26] ),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[0] ),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_fair_arb.i_lzc_lower.gen_lzc.in_tmp ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\i_snitch.i_snitch_regfile.mem[66] ),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\i_snitch.i_snitch_regfile.mem[354] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[35] ),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\rsp_data_q[10] ),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\i_snitch.i_snitch_regfile.mem[357] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\i_snitch.i_snitch_regfile.mem[228] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\i_snitch.i_snitch_regfile.mem[418] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\i_snitch.i_snitch_regfile.mem[37] ),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\i_snitch.i_snitch_regfile.mem[386] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[27] ),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\rsp_data_q[9] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\rsp_data_q[9]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\rsp_data_q[27] ),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\i_snitch.inst_addr_o[24] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\rsp_data_q[25] ),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\rsp_data_q[25]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\rsp_data_q[17] ),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\rsp_data_q[17]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\i_snitch.i_snitch_regfile.mem[299] ),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\i_snitch.i_snitch_regfile.mem[55] ),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\i_snitch.i_snitch_regfile.mem[101] ),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\rsp_data_q[0] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\i_snitch.inst_addr_o[18] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\i_snitch.i_snitch_regfile.mem[423] ),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold1325 (.A(\i_snitch.i_snitch_regfile.mem[226] ),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\i_snitch.i_snitch_regfile.mem[98] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\i_snitch.i_snitch_regfile.mem[259] ),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\i_snitch.i_snitch_regfile.mem[195] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\i_req_arb.data_i[41] ),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\rsp_data_q[19] ),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\i_snitch.inst_addr_o[14] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\i_snitch.i_snitch_regfile.mem[99] ),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\rsp_data_q[5] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\rsp_data_q[5]_sg13g2_dfrbpq_1_Q_D_sg13g2_inv_1_Y_A ),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\i_snitch.gpr_waddr[6] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\i_snitch.i_snitch_regfile.mem[229] ),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\rsp_data_q[2] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\i_snitch.i_snitch_regfile.mem[133] ),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\i_snitch.i_snitch_regfile.mem[403] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\i_snitch.inst_addr_o[23] ),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\i_snitch.inst_addr_o[26] ),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[30] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\i_snitch.inst_addr_o[13] ),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[6] ),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[15] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\i_req_arb.data_i[37] ),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\i_snitch.i_snitch_regfile.mem[36] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[5] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\rsp_data_q[3] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold1350 (.A(\rsp_data_q[1] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[23] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\rsp_data_q[21] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\i_snitch.inst_addr_o[11] ),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\i_snitch.inst_addr_o[29] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_data_q[38] ),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\rsp_data_q[13] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\i_snitch.gpr_waddr[7] ),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\i_snitch.inst_addr_o[30] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\i_req_register.spill_register_flushable_i.gen_spill_reg.a_full_q ),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.lock_d_sg13g2_nor2_1_Y_A ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\i_req_arb.data_i[39] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\i_snitch.inst_addr_o[20] ),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\i_snitch.inst_addr_o[16] ),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\i_snitch.inst_addr_o[15] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\i_req_arb.gen_arbiter.gen_int_rr.gen_lock.req_q[1] ),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\i_req_arb.gen_arbiter.req_d[1]_sg13g2_or2_1_X_A ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\i_req_arb.gen_arbiter.req_d[1] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\i_snitch.inst_addr_o[12] ),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\i_snitch.inst_addr_o[28] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\i_snitch.gpr_waddr[5] ),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\i_snitch.i_snitch_lsu.metadata_q[3] ),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\i_snitch.i_snitch_lsu.metadata_q[2] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\i_req_arb.data_i[43] ),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\i_snitch.inst_addr_o[22] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\i_snitch.i_snitch_lsu.handshake_pending_q ),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold1376 (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\i_inst_register.spill_register_flushable_i.gen_spill_reg.a_data_q[20] ),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold1378 (.A(data_pvalid_sg13g2_nor2_1_A_Y_sg13g2_dfrbpq_1_D_Q),
    .X(net1410));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_176 ();
 sg13g2_decap_8 FILLER_0_183 ();
 sg13g2_fill_1 FILLER_0_190 ();
 sg13g2_decap_8 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_decap_8 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_216 ();
 sg13g2_decap_8 FILLER_0_223 ();
 sg13g2_decap_8 FILLER_0_230 ();
 sg13g2_fill_1 FILLER_0_237 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_fill_2 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_fill_2 FILLER_0_292 ();
 sg13g2_fill_1 FILLER_0_294 ();
 sg13g2_fill_2 FILLER_0_303 ();
 sg13g2_fill_2 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_8 FILLER_0_351 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_365 ();
 sg13g2_decap_8 FILLER_0_372 ();
 sg13g2_decap_8 FILLER_0_379 ();
 sg13g2_decap_8 FILLER_0_386 ();
 sg13g2_decap_8 FILLER_0_393 ();
 sg13g2_decap_8 FILLER_0_400 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_8 FILLER_0_414 ();
 sg13g2_decap_4 FILLER_0_421 ();
 sg13g2_fill_2 FILLER_0_425 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_8 FILLER_0_468 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_fill_2 FILLER_0_482 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_fill_2 FILLER_0_539 ();
 sg13g2_fill_1 FILLER_0_541 ();
 sg13g2_decap_8 FILLER_0_569 ();
 sg13g2_decap_8 FILLER_0_576 ();
 sg13g2_decap_8 FILLER_0_583 ();
 sg13g2_decap_8 FILLER_0_590 ();
 sg13g2_decap_8 FILLER_0_597 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_8 FILLER_0_618 ();
 sg13g2_decap_8 FILLER_0_625 ();
 sg13g2_decap_8 FILLER_0_632 ();
 sg13g2_decap_8 FILLER_0_639 ();
 sg13g2_decap_8 FILLER_0_646 ();
 sg13g2_decap_8 FILLER_0_653 ();
 sg13g2_decap_8 FILLER_0_660 ();
 sg13g2_decap_8 FILLER_0_667 ();
 sg13g2_decap_8 FILLER_0_674 ();
 sg13g2_decap_8 FILLER_0_681 ();
 sg13g2_decap_8 FILLER_0_688 ();
 sg13g2_decap_8 FILLER_0_695 ();
 sg13g2_decap_8 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_709 ();
 sg13g2_decap_8 FILLER_0_716 ();
 sg13g2_decap_8 FILLER_0_723 ();
 sg13g2_decap_8 FILLER_0_730 ();
 sg13g2_decap_8 FILLER_0_737 ();
 sg13g2_decap_8 FILLER_0_744 ();
 sg13g2_decap_8 FILLER_0_751 ();
 sg13g2_decap_8 FILLER_0_758 ();
 sg13g2_decap_8 FILLER_0_765 ();
 sg13g2_decap_8 FILLER_0_772 ();
 sg13g2_decap_8 FILLER_0_779 ();
 sg13g2_decap_8 FILLER_0_786 ();
 sg13g2_decap_8 FILLER_0_793 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_decap_8 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_821 ();
 sg13g2_decap_8 FILLER_0_828 ();
 sg13g2_decap_8 FILLER_0_835 ();
 sg13g2_decap_8 FILLER_0_842 ();
 sg13g2_decap_8 FILLER_0_849 ();
 sg13g2_decap_8 FILLER_0_856 ();
 sg13g2_decap_8 FILLER_0_863 ();
 sg13g2_decap_8 FILLER_0_870 ();
 sg13g2_decap_8 FILLER_0_877 ();
 sg13g2_decap_8 FILLER_0_884 ();
 sg13g2_decap_8 FILLER_0_891 ();
 sg13g2_decap_8 FILLER_0_898 ();
 sg13g2_decap_8 FILLER_0_905 ();
 sg13g2_decap_8 FILLER_0_912 ();
 sg13g2_decap_8 FILLER_0_919 ();
 sg13g2_decap_8 FILLER_0_926 ();
 sg13g2_decap_8 FILLER_0_933 ();
 sg13g2_decap_8 FILLER_0_940 ();
 sg13g2_decap_8 FILLER_0_947 ();
 sg13g2_decap_8 FILLER_0_954 ();
 sg13g2_decap_8 FILLER_0_961 ();
 sg13g2_decap_8 FILLER_0_968 ();
 sg13g2_decap_8 FILLER_0_975 ();
 sg13g2_decap_8 FILLER_0_982 ();
 sg13g2_decap_8 FILLER_0_989 ();
 sg13g2_decap_8 FILLER_0_996 ();
 sg13g2_decap_8 FILLER_0_1003 ();
 sg13g2_decap_8 FILLER_0_1010 ();
 sg13g2_decap_8 FILLER_0_1017 ();
 sg13g2_decap_4 FILLER_0_1024 ();
 sg13g2_fill_1 FILLER_0_1028 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_4 FILLER_1_147 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_2 FILLER_1_261 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_fill_2 FILLER_1_295 ();
 sg13g2_fill_1 FILLER_1_297 ();
 sg13g2_decap_4 FILLER_1_415 ();
 sg13g2_fill_1 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_1_460 ();
 sg13g2_fill_2 FILLER_1_467 ();
 sg13g2_fill_1 FILLER_1_469 ();
 sg13g2_fill_2 FILLER_1_555 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_8 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_580 ();
 sg13g2_decap_8 FILLER_1_587 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_8 FILLER_1_601 ();
 sg13g2_decap_8 FILLER_1_608 ();
 sg13g2_decap_8 FILLER_1_615 ();
 sg13g2_decap_8 FILLER_1_622 ();
 sg13g2_decap_8 FILLER_1_629 ();
 sg13g2_decap_8 FILLER_1_636 ();
 sg13g2_decap_8 FILLER_1_643 ();
 sg13g2_decap_8 FILLER_1_650 ();
 sg13g2_decap_8 FILLER_1_657 ();
 sg13g2_decap_8 FILLER_1_664 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_decap_8 FILLER_1_685 ();
 sg13g2_decap_8 FILLER_1_692 ();
 sg13g2_decap_8 FILLER_1_699 ();
 sg13g2_decap_8 FILLER_1_706 ();
 sg13g2_decap_8 FILLER_1_713 ();
 sg13g2_decap_8 FILLER_1_720 ();
 sg13g2_decap_8 FILLER_1_727 ();
 sg13g2_decap_8 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_741 ();
 sg13g2_decap_8 FILLER_1_748 ();
 sg13g2_decap_8 FILLER_1_755 ();
 sg13g2_decap_8 FILLER_1_762 ();
 sg13g2_decap_8 FILLER_1_769 ();
 sg13g2_decap_8 FILLER_1_776 ();
 sg13g2_decap_8 FILLER_1_783 ();
 sg13g2_decap_8 FILLER_1_790 ();
 sg13g2_decap_8 FILLER_1_797 ();
 sg13g2_decap_8 FILLER_1_804 ();
 sg13g2_decap_8 FILLER_1_811 ();
 sg13g2_decap_8 FILLER_1_818 ();
 sg13g2_decap_8 FILLER_1_825 ();
 sg13g2_decap_8 FILLER_1_832 ();
 sg13g2_decap_8 FILLER_1_839 ();
 sg13g2_decap_8 FILLER_1_846 ();
 sg13g2_decap_8 FILLER_1_853 ();
 sg13g2_decap_8 FILLER_1_860 ();
 sg13g2_decap_8 FILLER_1_867 ();
 sg13g2_decap_8 FILLER_1_874 ();
 sg13g2_decap_8 FILLER_1_881 ();
 sg13g2_decap_8 FILLER_1_888 ();
 sg13g2_decap_8 FILLER_1_895 ();
 sg13g2_decap_8 FILLER_1_902 ();
 sg13g2_decap_8 FILLER_1_909 ();
 sg13g2_decap_8 FILLER_1_916 ();
 sg13g2_decap_8 FILLER_1_923 ();
 sg13g2_decap_8 FILLER_1_930 ();
 sg13g2_decap_8 FILLER_1_937 ();
 sg13g2_decap_8 FILLER_1_944 ();
 sg13g2_decap_8 FILLER_1_951 ();
 sg13g2_decap_8 FILLER_1_958 ();
 sg13g2_decap_8 FILLER_1_965 ();
 sg13g2_decap_8 FILLER_1_972 ();
 sg13g2_decap_8 FILLER_1_979 ();
 sg13g2_decap_8 FILLER_1_986 ();
 sg13g2_decap_8 FILLER_1_993 ();
 sg13g2_decap_8 FILLER_1_1000 ();
 sg13g2_decap_8 FILLER_1_1007 ();
 sg13g2_decap_8 FILLER_1_1014 ();
 sg13g2_decap_8 FILLER_1_1021 ();
 sg13g2_fill_1 FILLER_1_1028 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_4 FILLER_2_137 ();
 sg13g2_fill_1 FILLER_2_141 ();
 sg13g2_fill_1 FILLER_2_169 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_232 ();
 sg13g2_fill_2 FILLER_2_246 ();
 sg13g2_fill_2 FILLER_2_306 ();
 sg13g2_fill_1 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_348 ();
 sg13g2_fill_2 FILLER_2_355 ();
 sg13g2_fill_1 FILLER_2_384 ();
 sg13g2_fill_1 FILLER_2_418 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_4 FILLER_2_460 ();
 sg13g2_fill_2 FILLER_2_464 ();
 sg13g2_fill_1 FILLER_2_480 ();
 sg13g2_fill_2 FILLER_2_496 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_fill_1 FILLER_2_527 ();
 sg13g2_fill_1 FILLER_2_577 ();
 sg13g2_decap_8 FILLER_2_582 ();
 sg13g2_decap_8 FILLER_2_589 ();
 sg13g2_decap_8 FILLER_2_600 ();
 sg13g2_decap_8 FILLER_2_607 ();
 sg13g2_decap_8 FILLER_2_614 ();
 sg13g2_decap_8 FILLER_2_621 ();
 sg13g2_decap_8 FILLER_2_628 ();
 sg13g2_decap_8 FILLER_2_635 ();
 sg13g2_decap_8 FILLER_2_642 ();
 sg13g2_decap_8 FILLER_2_649 ();
 sg13g2_decap_8 FILLER_2_656 ();
 sg13g2_decap_8 FILLER_2_663 ();
 sg13g2_decap_8 FILLER_2_670 ();
 sg13g2_decap_8 FILLER_2_677 ();
 sg13g2_decap_8 FILLER_2_684 ();
 sg13g2_decap_8 FILLER_2_691 ();
 sg13g2_decap_8 FILLER_2_698 ();
 sg13g2_decap_8 FILLER_2_705 ();
 sg13g2_decap_8 FILLER_2_712 ();
 sg13g2_decap_8 FILLER_2_719 ();
 sg13g2_decap_4 FILLER_2_726 ();
 sg13g2_fill_2 FILLER_2_730 ();
 sg13g2_decap_8 FILLER_2_740 ();
 sg13g2_decap_8 FILLER_2_747 ();
 sg13g2_decap_8 FILLER_2_754 ();
 sg13g2_decap_8 FILLER_2_761 ();
 sg13g2_decap_8 FILLER_2_768 ();
 sg13g2_decap_8 FILLER_2_775 ();
 sg13g2_decap_8 FILLER_2_782 ();
 sg13g2_fill_2 FILLER_2_789 ();
 sg13g2_fill_1 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_796 ();
 sg13g2_decap_8 FILLER_2_803 ();
 sg13g2_decap_8 FILLER_2_810 ();
 sg13g2_decap_8 FILLER_2_817 ();
 sg13g2_decap_8 FILLER_2_824 ();
 sg13g2_decap_8 FILLER_2_831 ();
 sg13g2_decap_8 FILLER_2_838 ();
 sg13g2_decap_8 FILLER_2_845 ();
 sg13g2_decap_8 FILLER_2_852 ();
 sg13g2_decap_8 FILLER_2_859 ();
 sg13g2_decap_8 FILLER_2_866 ();
 sg13g2_decap_8 FILLER_2_873 ();
 sg13g2_decap_8 FILLER_2_880 ();
 sg13g2_decap_8 FILLER_2_887 ();
 sg13g2_decap_8 FILLER_2_894 ();
 sg13g2_decap_8 FILLER_2_901 ();
 sg13g2_decap_8 FILLER_2_908 ();
 sg13g2_decap_8 FILLER_2_915 ();
 sg13g2_decap_8 FILLER_2_922 ();
 sg13g2_decap_8 FILLER_2_929 ();
 sg13g2_decap_8 FILLER_2_936 ();
 sg13g2_decap_8 FILLER_2_943 ();
 sg13g2_decap_8 FILLER_2_950 ();
 sg13g2_decap_8 FILLER_2_957 ();
 sg13g2_decap_8 FILLER_2_964 ();
 sg13g2_decap_8 FILLER_2_971 ();
 sg13g2_decap_8 FILLER_2_978 ();
 sg13g2_decap_8 FILLER_2_985 ();
 sg13g2_decap_8 FILLER_2_992 ();
 sg13g2_decap_8 FILLER_2_999 ();
 sg13g2_decap_8 FILLER_2_1006 ();
 sg13g2_decap_8 FILLER_2_1013 ();
 sg13g2_decap_8 FILLER_2_1020 ();
 sg13g2_fill_2 FILLER_2_1027 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_167 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_fill_2 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_225 ();
 sg13g2_decap_8 FILLER_3_236 ();
 sg13g2_fill_1 FILLER_3_243 ();
 sg13g2_fill_2 FILLER_3_252 ();
 sg13g2_fill_2 FILLER_3_258 ();
 sg13g2_fill_2 FILLER_3_276 ();
 sg13g2_fill_1 FILLER_3_278 ();
 sg13g2_fill_1 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_314 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_decap_4 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_369 ();
 sg13g2_fill_2 FILLER_3_383 ();
 sg13g2_fill_1 FILLER_3_385 ();
 sg13g2_fill_1 FILLER_3_422 ();
 sg13g2_decap_4 FILLER_3_433 ();
 sg13g2_fill_2 FILLER_3_437 ();
 sg13g2_decap_8 FILLER_3_460 ();
 sg13g2_fill_2 FILLER_3_467 ();
 sg13g2_fill_2 FILLER_3_486 ();
 sg13g2_decap_8 FILLER_3_492 ();
 sg13g2_fill_2 FILLER_3_499 ();
 sg13g2_fill_1 FILLER_3_575 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_646 ();
 sg13g2_decap_8 FILLER_3_653 ();
 sg13g2_decap_8 FILLER_3_660 ();
 sg13g2_decap_8 FILLER_3_667 ();
 sg13g2_decap_8 FILLER_3_674 ();
 sg13g2_decap_4 FILLER_3_681 ();
 sg13g2_fill_2 FILLER_3_685 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_fill_2 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_758 ();
 sg13g2_decap_8 FILLER_3_765 ();
 sg13g2_decap_8 FILLER_3_772 ();
 sg13g2_decap_4 FILLER_3_779 ();
 sg13g2_fill_1 FILLER_3_783 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_8 FILLER_3_913 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_decap_8 FILLER_3_927 ();
 sg13g2_decap_8 FILLER_3_934 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_8 FILLER_3_976 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_219 ();
 sg13g2_decap_4 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_268 ();
 sg13g2_decap_8 FILLER_4_283 ();
 sg13g2_decap_8 FILLER_4_290 ();
 sg13g2_decap_4 FILLER_4_297 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_4 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_4 FILLER_4_357 ();
 sg13g2_fill_2 FILLER_4_361 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_2 FILLER_4_396 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_fill_1 FILLER_4_473 ();
 sg13g2_fill_2 FILLER_4_537 ();
 sg13g2_fill_2 FILLER_4_578 ();
 sg13g2_fill_1 FILLER_4_580 ();
 sg13g2_fill_2 FILLER_4_617 ();
 sg13g2_fill_1 FILLER_4_619 ();
 sg13g2_decap_8 FILLER_4_647 ();
 sg13g2_decap_8 FILLER_4_654 ();
 sg13g2_decap_8 FILLER_4_661 ();
 sg13g2_decap_8 FILLER_4_668 ();
 sg13g2_decap_8 FILLER_4_675 ();
 sg13g2_fill_2 FILLER_4_682 ();
 sg13g2_fill_1 FILLER_4_697 ();
 sg13g2_fill_1 FILLER_4_725 ();
 sg13g2_fill_2 FILLER_4_741 ();
 sg13g2_fill_1 FILLER_4_743 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_4 FILLER_4_884 ();
 sg13g2_fill_1 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_920 ();
 sg13g2_decap_8 FILLER_4_927 ();
 sg13g2_decap_8 FILLER_4_934 ();
 sg13g2_decap_8 FILLER_4_941 ();
 sg13g2_decap_8 FILLER_4_948 ();
 sg13g2_decap_8 FILLER_4_955 ();
 sg13g2_decap_8 FILLER_4_962 ();
 sg13g2_decap_8 FILLER_4_969 ();
 sg13g2_decap_8 FILLER_4_976 ();
 sg13g2_decap_8 FILLER_4_983 ();
 sg13g2_decap_8 FILLER_4_990 ();
 sg13g2_decap_8 FILLER_4_997 ();
 sg13g2_decap_8 FILLER_4_1004 ();
 sg13g2_decap_8 FILLER_4_1011 ();
 sg13g2_decap_8 FILLER_4_1018 ();
 sg13g2_decap_4 FILLER_4_1025 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_4 FILLER_5_158 ();
 sg13g2_fill_2 FILLER_5_162 ();
 sg13g2_decap_4 FILLER_5_178 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_5_203 ();
 sg13g2_decap_4 FILLER_5_209 ();
 sg13g2_fill_2 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_242 ();
 sg13g2_fill_1 FILLER_5_244 ();
 sg13g2_fill_2 FILLER_5_258 ();
 sg13g2_fill_1 FILLER_5_275 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_4 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_436 ();
 sg13g2_fill_2 FILLER_5_470 ();
 sg13g2_fill_1 FILLER_5_472 ();
 sg13g2_fill_2 FILLER_5_479 ();
 sg13g2_fill_1 FILLER_5_481 ();
 sg13g2_fill_1 FILLER_5_495 ();
 sg13g2_fill_2 FILLER_5_534 ();
 sg13g2_fill_2 FILLER_5_542 ();
 sg13g2_fill_2 FILLER_5_583 ();
 sg13g2_fill_2 FILLER_5_621 ();
 sg13g2_decap_8 FILLER_5_642 ();
 sg13g2_fill_1 FILLER_5_649 ();
 sg13g2_fill_1 FILLER_5_663 ();
 sg13g2_fill_2 FILLER_5_691 ();
 sg13g2_fill_1 FILLER_5_693 ();
 sg13g2_fill_2 FILLER_5_721 ();
 sg13g2_fill_2 FILLER_5_789 ();
 sg13g2_fill_1 FILLER_5_791 ();
 sg13g2_fill_1 FILLER_5_870 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_167 ();
 sg13g2_fill_2 FILLER_6_214 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_258 ();
 sg13g2_fill_1 FILLER_6_260 ();
 sg13g2_decap_4 FILLER_6_301 ();
 sg13g2_decap_4 FILLER_6_356 ();
 sg13g2_fill_1 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_370 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_4 FILLER_6_387 ();
 sg13g2_fill_1 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_6_412 ();
 sg13g2_fill_2 FILLER_6_419 ();
 sg13g2_fill_1 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_fill_1 FILLER_6_430 ();
 sg13g2_decap_4 FILLER_6_458 ();
 sg13g2_fill_2 FILLER_6_471 ();
 sg13g2_fill_2 FILLER_6_481 ();
 sg13g2_fill_1 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_503 ();
 sg13g2_fill_2 FILLER_6_510 ();
 sg13g2_fill_1 FILLER_6_533 ();
 sg13g2_fill_1 FILLER_6_538 ();
 sg13g2_fill_2 FILLER_6_570 ();
 sg13g2_fill_1 FILLER_6_572 ();
 sg13g2_decap_8 FILLER_6_604 ();
 sg13g2_decap_4 FILLER_6_611 ();
 sg13g2_fill_1 FILLER_6_615 ();
 sg13g2_decap_4 FILLER_6_624 ();
 sg13g2_fill_1 FILLER_6_628 ();
 sg13g2_fill_2 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_644 ();
 sg13g2_decap_4 FILLER_6_676 ();
 sg13g2_fill_1 FILLER_6_680 ();
 sg13g2_decap_8 FILLER_6_685 ();
 sg13g2_decap_8 FILLER_6_692 ();
 sg13g2_decap_8 FILLER_6_699 ();
 sg13g2_fill_2 FILLER_6_706 ();
 sg13g2_fill_2 FILLER_6_725 ();
 sg13g2_fill_1 FILLER_6_727 ();
 sg13g2_fill_1 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_758 ();
 sg13g2_decap_4 FILLER_6_765 ();
 sg13g2_fill_1 FILLER_6_782 ();
 sg13g2_fill_2 FILLER_6_817 ();
 sg13g2_fill_2 FILLER_6_872 ();
 sg13g2_fill_1 FILLER_6_874 ();
 sg13g2_fill_2 FILLER_6_885 ();
 sg13g2_fill_1 FILLER_6_887 ();
 sg13g2_fill_2 FILLER_6_903 ();
 sg13g2_fill_1 FILLER_6_905 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_4 ();
 sg13g2_decap_8 FILLER_7_11 ();
 sg13g2_decap_8 FILLER_7_18 ();
 sg13g2_decap_8 FILLER_7_25 ();
 sg13g2_decap_8 FILLER_7_32 ();
 sg13g2_decap_8 FILLER_7_39 ();
 sg13g2_decap_8 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_67 ();
 sg13g2_fill_2 FILLER_7_74 ();
 sg13g2_fill_2 FILLER_7_94 ();
 sg13g2_decap_8 FILLER_7_108 ();
 sg13g2_decap_4 FILLER_7_115 ();
 sg13g2_decap_8 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_137 ();
 sg13g2_decap_4 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_220 ();
 sg13g2_fill_1 FILLER_7_222 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_4 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_277 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_fill_2 FILLER_7_294 ();
 sg13g2_decap_4 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_4 FILLER_7_322 ();
 sg13g2_fill_1 FILLER_7_329 ();
 sg13g2_decap_4 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_fill_2 FILLER_7_411 ();
 sg13g2_fill_1 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_433 ();
 sg13g2_decap_4 FILLER_7_445 ();
 sg13g2_fill_1 FILLER_7_449 ();
 sg13g2_fill_2 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_460 ();
 sg13g2_decap_8 FILLER_7_467 ();
 sg13g2_decap_4 FILLER_7_474 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_fill_1 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_568 ();
 sg13g2_decap_8 FILLER_7_575 ();
 sg13g2_decap_4 FILLER_7_582 ();
 sg13g2_decap_4 FILLER_7_592 ();
 sg13g2_fill_1 FILLER_7_596 ();
 sg13g2_fill_1 FILLER_7_619 ();
 sg13g2_decap_8 FILLER_7_633 ();
 sg13g2_fill_1 FILLER_7_640 ();
 sg13g2_fill_2 FILLER_7_658 ();
 sg13g2_fill_2 FILLER_7_673 ();
 sg13g2_fill_1 FILLER_7_675 ();
 sg13g2_fill_2 FILLER_7_682 ();
 sg13g2_fill_1 FILLER_7_684 ();
 sg13g2_decap_4 FILLER_7_694 ();
 sg13g2_fill_2 FILLER_7_711 ();
 sg13g2_decap_4 FILLER_7_745 ();
 sg13g2_decap_8 FILLER_7_753 ();
 sg13g2_decap_8 FILLER_7_760 ();
 sg13g2_decap_8 FILLER_7_767 ();
 sg13g2_fill_2 FILLER_7_774 ();
 sg13g2_fill_1 FILLER_7_776 ();
 sg13g2_decap_8 FILLER_7_797 ();
 sg13g2_decap_4 FILLER_7_808 ();
 sg13g2_decap_8 FILLER_7_822 ();
 sg13g2_fill_2 FILLER_7_846 ();
 sg13g2_fill_1 FILLER_7_848 ();
 sg13g2_decap_4 FILLER_7_855 ();
 sg13g2_fill_2 FILLER_7_859 ();
 sg13g2_fill_1 FILLER_7_870 ();
 sg13g2_fill_2 FILLER_7_892 ();
 sg13g2_fill_1 FILLER_7_894 ();
 sg13g2_fill_1 FILLER_7_899 ();
 sg13g2_fill_1 FILLER_7_908 ();
 sg13g2_fill_1 FILLER_7_948 ();
 sg13g2_decap_8 FILLER_7_976 ();
 sg13g2_decap_8 FILLER_7_983 ();
 sg13g2_decap_8 FILLER_7_990 ();
 sg13g2_decap_8 FILLER_7_997 ();
 sg13g2_decap_8 FILLER_7_1004 ();
 sg13g2_decap_8 FILLER_7_1011 ();
 sg13g2_decap_8 FILLER_7_1018 ();
 sg13g2_decap_4 FILLER_7_1025 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_fill_2 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_65 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_135 ();
 sg13g2_decap_8 FILLER_8_142 ();
 sg13g2_decap_8 FILLER_8_149 ();
 sg13g2_decap_8 FILLER_8_156 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_2 FILLER_8_213 ();
 sg13g2_fill_1 FILLER_8_248 ();
 sg13g2_decap_4 FILLER_8_274 ();
 sg13g2_fill_2 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_307 ();
 sg13g2_fill_2 FILLER_8_313 ();
 sg13g2_fill_1 FILLER_8_315 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_398 ();
 sg13g2_fill_1 FILLER_8_426 ();
 sg13g2_fill_1 FILLER_8_448 ();
 sg13g2_fill_2 FILLER_8_466 ();
 sg13g2_decap_4 FILLER_8_503 ();
 sg13g2_fill_2 FILLER_8_507 ();
 sg13g2_decap_4 FILLER_8_512 ();
 sg13g2_decap_8 FILLER_8_540 ();
 sg13g2_fill_2 FILLER_8_547 ();
 sg13g2_fill_1 FILLER_8_549 ();
 sg13g2_decap_4 FILLER_8_554 ();
 sg13g2_fill_1 FILLER_8_558 ();
 sg13g2_decap_4 FILLER_8_568 ();
 sg13g2_fill_2 FILLER_8_585 ();
 sg13g2_decap_4 FILLER_8_600 ();
 sg13g2_fill_1 FILLER_8_608 ();
 sg13g2_decap_8 FILLER_8_659 ();
 sg13g2_decap_4 FILLER_8_666 ();
 sg13g2_fill_2 FILLER_8_680 ();
 sg13g2_fill_2 FILLER_8_709 ();
 sg13g2_fill_2 FILLER_8_742 ();
 sg13g2_fill_1 FILLER_8_744 ();
 sg13g2_fill_2 FILLER_8_776 ();
 sg13g2_fill_1 FILLER_8_778 ();
 sg13g2_fill_2 FILLER_8_815 ();
 sg13g2_fill_1 FILLER_8_817 ();
 sg13g2_decap_8 FILLER_8_845 ();
 sg13g2_fill_2 FILLER_8_852 ();
 sg13g2_fill_2 FILLER_8_907 ();
 sg13g2_fill_1 FILLER_8_909 ();
 sg13g2_fill_2 FILLER_8_940 ();
 sg13g2_decap_8 FILLER_8_969 ();
 sg13g2_decap_8 FILLER_8_976 ();
 sg13g2_decap_8 FILLER_8_983 ();
 sg13g2_decap_8 FILLER_8_990 ();
 sg13g2_decap_8 FILLER_8_997 ();
 sg13g2_decap_8 FILLER_8_1004 ();
 sg13g2_decap_8 FILLER_8_1011 ();
 sg13g2_decap_8 FILLER_8_1018 ();
 sg13g2_decap_4 FILLER_8_1025 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_4 FILLER_9_49 ();
 sg13g2_fill_2 FILLER_9_80 ();
 sg13g2_decap_8 FILLER_9_128 ();
 sg13g2_decap_4 FILLER_9_135 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_222 ();
 sg13g2_fill_2 FILLER_9_241 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_297 ();
 sg13g2_fill_1 FILLER_9_326 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_fill_2 FILLER_9_405 ();
 sg13g2_decap_4 FILLER_9_411 ();
 sg13g2_fill_2 FILLER_9_415 ();
 sg13g2_fill_2 FILLER_9_432 ();
 sg13g2_decap_4 FILLER_9_443 ();
 sg13g2_fill_1 FILLER_9_447 ();
 sg13g2_fill_2 FILLER_9_453 ();
 sg13g2_fill_1 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_4 FILLER_9_483 ();
 sg13g2_fill_1 FILLER_9_487 ();
 sg13g2_fill_2 FILLER_9_494 ();
 sg13g2_fill_1 FILLER_9_496 ();
 sg13g2_decap_8 FILLER_9_506 ();
 sg13g2_decap_4 FILLER_9_513 ();
 sg13g2_fill_1 FILLER_9_517 ();
 sg13g2_fill_1 FILLER_9_544 ();
 sg13g2_decap_8 FILLER_9_572 ();
 sg13g2_decap_4 FILLER_9_579 ();
 sg13g2_fill_2 FILLER_9_583 ();
 sg13g2_fill_1 FILLER_9_604 ();
 sg13g2_fill_2 FILLER_9_624 ();
 sg13g2_decap_4 FILLER_9_635 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_fill_2 FILLER_9_700 ();
 sg13g2_fill_1 FILLER_9_702 ();
 sg13g2_decap_8 FILLER_9_720 ();
 sg13g2_decap_8 FILLER_9_727 ();
 sg13g2_decap_8 FILLER_9_734 ();
 sg13g2_fill_2 FILLER_9_741 ();
 sg13g2_fill_1 FILLER_9_747 ();
 sg13g2_decap_8 FILLER_9_754 ();
 sg13g2_fill_2 FILLER_9_761 ();
 sg13g2_decap_8 FILLER_9_772 ();
 sg13g2_decap_4 FILLER_9_779 ();
 sg13g2_decap_8 FILLER_9_787 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_fill_2 FILLER_9_839 ();
 sg13g2_fill_1 FILLER_9_841 ();
 sg13g2_decap_8 FILLER_9_873 ();
 sg13g2_decap_4 FILLER_9_880 ();
 sg13g2_fill_1 FILLER_9_968 ();
 sg13g2_decap_8 FILLER_9_978 ();
 sg13g2_decap_8 FILLER_9_985 ();
 sg13g2_decap_8 FILLER_9_992 ();
 sg13g2_decap_8 FILLER_9_999 ();
 sg13g2_decap_8 FILLER_9_1006 ();
 sg13g2_decap_8 FILLER_9_1013 ();
 sg13g2_decap_8 FILLER_9_1020 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_fill_2 FILLER_10_25 ();
 sg13g2_fill_2 FILLER_10_54 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_2 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_fill_1 FILLER_10_115 ();
 sg13g2_decap_8 FILLER_10_152 ();
 sg13g2_fill_1 FILLER_10_159 ();
 sg13g2_decap_8 FILLER_10_204 ();
 sg13g2_decap_8 FILLER_10_211 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_250 ();
 sg13g2_fill_1 FILLER_10_252 ();
 sg13g2_decap_4 FILLER_10_281 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_289 ();
 sg13g2_decap_4 FILLER_10_295 ();
 sg13g2_fill_1 FILLER_10_299 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_decap_4 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_4 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_4 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_4 FILLER_10_386 ();
 sg13g2_fill_2 FILLER_10_390 ();
 sg13g2_fill_1 FILLER_10_405 ();
 sg13g2_fill_1 FILLER_10_419 ();
 sg13g2_fill_2 FILLER_10_424 ();
 sg13g2_fill_1 FILLER_10_426 ();
 sg13g2_fill_2 FILLER_10_440 ();
 sg13g2_fill_1 FILLER_10_442 ();
 sg13g2_fill_2 FILLER_10_453 ();
 sg13g2_decap_4 FILLER_10_464 ();
 sg13g2_fill_1 FILLER_10_491 ();
 sg13g2_fill_1 FILLER_10_501 ();
 sg13g2_decap_4 FILLER_10_506 ();
 sg13g2_fill_1 FILLER_10_533 ();
 sg13g2_fill_1 FILLER_10_540 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_fill_2 FILLER_10_594 ();
 sg13g2_fill_2 FILLER_10_623 ();
 sg13g2_fill_1 FILLER_10_625 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_fill_2 FILLER_10_637 ();
 sg13g2_fill_1 FILLER_10_639 ();
 sg13g2_decap_4 FILLER_10_675 ();
 sg13g2_fill_1 FILLER_10_679 ();
 sg13g2_decap_4 FILLER_10_693 ();
 sg13g2_fill_1 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_fill_2 FILLER_10_732 ();
 sg13g2_fill_1 FILLER_10_734 ();
 sg13g2_decap_4 FILLER_10_766 ();
 sg13g2_decap_8 FILLER_10_797 ();
 sg13g2_decap_4 FILLER_10_804 ();
 sg13g2_fill_2 FILLER_10_845 ();
 sg13g2_fill_1 FILLER_10_847 ();
 sg13g2_decap_4 FILLER_10_858 ();
 sg13g2_decap_4 FILLER_10_871 ();
 sg13g2_decap_8 FILLER_10_878 ();
 sg13g2_fill_1 FILLER_10_885 ();
 sg13g2_fill_1 FILLER_10_932 ();
 sg13g2_fill_2 FILLER_10_948 ();
 sg13g2_fill_1 FILLER_10_967 ();
 sg13g2_decap_8 FILLER_10_999 ();
 sg13g2_decap_8 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1013 ();
 sg13g2_decap_8 FILLER_10_1020 ();
 sg13g2_fill_2 FILLER_10_1027 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_30 ();
 sg13g2_fill_1 FILLER_11_72 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_fill_1 FILLER_11_120 ();
 sg13g2_decap_8 FILLER_11_143 ();
 sg13g2_decap_8 FILLER_11_150 ();
 sg13g2_decap_4 FILLER_11_157 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_271 ();
 sg13g2_fill_1 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_4 FILLER_11_336 ();
 sg13g2_fill_1 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_fill_2 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_468 ();
 sg13g2_decap_8 FILLER_11_524 ();
 sg13g2_decap_8 FILLER_11_531 ();
 sg13g2_fill_2 FILLER_11_555 ();
 sg13g2_fill_2 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_607 ();
 sg13g2_fill_2 FILLER_11_614 ();
 sg13g2_fill_1 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_4 FILLER_11_651 ();
 sg13g2_fill_2 FILLER_11_772 ();
 sg13g2_fill_2 FILLER_11_778 ();
 sg13g2_fill_2 FILLER_11_816 ();
 sg13g2_fill_2 FILLER_11_850 ();
 sg13g2_fill_1 FILLER_11_852 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_fill_2 FILLER_11_954 ();
 sg13g2_fill_1 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_fill_1 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_8 ();
 sg13g2_fill_2 FILLER_12_15 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_112 ();
 sg13g2_fill_1 FILLER_12_114 ();
 sg13g2_decap_4 FILLER_12_147 ();
 sg13g2_fill_1 FILLER_12_151 ();
 sg13g2_fill_1 FILLER_12_213 ();
 sg13g2_decap_4 FILLER_12_232 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_decap_4 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_286 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_fill_2 FILLER_12_370 ();
 sg13g2_fill_1 FILLER_12_372 ();
 sg13g2_decap_4 FILLER_12_377 ();
 sg13g2_fill_2 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_fill_1 FILLER_12_421 ();
 sg13g2_decap_8 FILLER_12_439 ();
 sg13g2_decap_4 FILLER_12_459 ();
 sg13g2_fill_1 FILLER_12_475 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_526 ();
 sg13g2_fill_1 FILLER_12_579 ();
 sg13g2_fill_2 FILLER_12_603 ();
 sg13g2_fill_1 FILLER_12_605 ();
 sg13g2_fill_1 FILLER_12_632 ();
 sg13g2_fill_1 FILLER_12_639 ();
 sg13g2_fill_2 FILLER_12_653 ();
 sg13g2_decap_8 FILLER_12_671 ();
 sg13g2_fill_1 FILLER_12_678 ();
 sg13g2_fill_1 FILLER_12_692 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_fill_1 FILLER_12_756 ();
 sg13g2_decap_4 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_808 ();
 sg13g2_fill_1 FILLER_12_815 ();
 sg13g2_decap_4 FILLER_12_820 ();
 sg13g2_fill_2 FILLER_12_837 ();
 sg13g2_fill_1 FILLER_12_839 ();
 sg13g2_decap_4 FILLER_12_873 ();
 sg13g2_fill_1 FILLER_12_877 ();
 sg13g2_decap_4 FILLER_12_891 ();
 sg13g2_fill_1 FILLER_12_965 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_4 FILLER_12_984 ();
 sg13g2_fill_1 FILLER_12_988 ();
 sg13g2_fill_2 FILLER_12_1002 ();
 sg13g2_decap_8 FILLER_12_1013 ();
 sg13g2_decap_8 FILLER_12_1020 ();
 sg13g2_fill_2 FILLER_12_1027 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_39 ();
 sg13g2_fill_2 FILLER_13_43 ();
 sg13g2_decap_4 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_fill_1 FILLER_13_260 ();
 sg13g2_decap_8 FILLER_13_282 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_decap_4 FILLER_13_328 ();
 sg13g2_decap_8 FILLER_13_337 ();
 sg13g2_fill_2 FILLER_13_348 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_4 FILLER_13_384 ();
 sg13g2_decap_4 FILLER_13_412 ();
 sg13g2_fill_2 FILLER_13_416 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_4 FILLER_13_445 ();
 sg13g2_fill_1 FILLER_13_449 ();
 sg13g2_decap_4 FILLER_13_470 ();
 sg13g2_decap_8 FILLER_13_491 ();
 sg13g2_decap_4 FILLER_13_498 ();
 sg13g2_fill_1 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_fill_2 FILLER_13_573 ();
 sg13g2_fill_2 FILLER_13_598 ();
 sg13g2_fill_2 FILLER_13_618 ();
 sg13g2_fill_2 FILLER_13_654 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_fill_2 FILLER_13_693 ();
 sg13g2_decap_4 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_4 FILLER_13_833 ();
 sg13g2_fill_1 FILLER_13_850 ();
 sg13g2_fill_2 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_fill_2 FILLER_13_900 ();
 sg13g2_fill_1 FILLER_13_902 ();
 sg13g2_decap_8 FILLER_13_913 ();
 sg13g2_fill_2 FILLER_13_929 ();
 sg13g2_fill_1 FILLER_13_931 ();
 sg13g2_decap_8 FILLER_13_953 ();
 sg13g2_decap_8 FILLER_13_960 ();
 sg13g2_decap_8 FILLER_13_967 ();
 sg13g2_decap_8 FILLER_13_1013 ();
 sg13g2_decap_8 FILLER_13_1020 ();
 sg13g2_fill_2 FILLER_13_1027 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_29 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_1 FILLER_14_124 ();
 sg13g2_fill_2 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_155 ();
 sg13g2_decap_8 FILLER_14_162 ();
 sg13g2_fill_2 FILLER_14_186 ();
 sg13g2_fill_1 FILLER_14_188 ();
 sg13g2_decap_8 FILLER_14_262 ();
 sg13g2_fill_1 FILLER_14_273 ();
 sg13g2_decap_4 FILLER_14_280 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_decap_4 FILLER_14_326 ();
 sg13g2_fill_1 FILLER_14_351 ();
 sg13g2_decap_8 FILLER_14_365 ();
 sg13g2_decap_4 FILLER_14_372 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_415 ();
 sg13g2_decap_8 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_14_433 ();
 sg13g2_fill_1 FILLER_14_440 ();
 sg13g2_fill_2 FILLER_14_445 ();
 sg13g2_fill_1 FILLER_14_447 ();
 sg13g2_fill_1 FILLER_14_454 ();
 sg13g2_fill_2 FILLER_14_468 ();
 sg13g2_fill_1 FILLER_14_497 ();
 sg13g2_fill_2 FILLER_14_511 ();
 sg13g2_fill_1 FILLER_14_513 ();
 sg13g2_decap_4 FILLER_14_533 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_fill_1 FILLER_14_552 ();
 sg13g2_fill_2 FILLER_14_591 ();
 sg13g2_fill_1 FILLER_14_593 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_4 FILLER_14_664 ();
 sg13g2_fill_2 FILLER_14_705 ();
 sg13g2_fill_1 FILLER_14_707 ();
 sg13g2_fill_1 FILLER_14_733 ();
 sg13g2_fill_1 FILLER_14_744 ();
 sg13g2_decap_4 FILLER_14_762 ();
 sg13g2_decap_8 FILLER_14_772 ();
 sg13g2_fill_2 FILLER_14_779 ();
 sg13g2_fill_1 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_4 FILLER_14_798 ();
 sg13g2_fill_1 FILLER_14_802 ();
 sg13g2_fill_2 FILLER_14_809 ();
 sg13g2_fill_2 FILLER_14_851 ();
 sg13g2_fill_2 FILLER_14_889 ();
 sg13g2_fill_1 FILLER_14_891 ();
 sg13g2_decap_8 FILLER_14_905 ();
 sg13g2_decap_8 FILLER_14_912 ();
 sg13g2_fill_2 FILLER_14_919 ();
 sg13g2_fill_1 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_fill_2 FILLER_14_935 ();
 sg13g2_fill_1 FILLER_14_967 ();
 sg13g2_fill_1 FILLER_14_974 ();
 sg13g2_fill_1 FILLER_14_983 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_2 ();
 sg13g2_fill_2 FILLER_15_22 ();
 sg13g2_fill_1 FILLER_15_24 ();
 sg13g2_fill_2 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_67 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_129 ();
 sg13g2_decap_4 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_181 ();
 sg13g2_decap_8 FILLER_15_188 ();
 sg13g2_decap_8 FILLER_15_195 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_4 FILLER_15_218 ();
 sg13g2_fill_2 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_241 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_4 FILLER_15_255 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_300 ();
 sg13g2_decap_4 FILLER_15_316 ();
 sg13g2_fill_2 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_331 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_352 ();
 sg13g2_decap_8 FILLER_15_380 ();
 sg13g2_decap_4 FILLER_15_387 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_fill_1 FILLER_15_402 ();
 sg13g2_fill_1 FILLER_15_430 ();
 sg13g2_decap_8 FILLER_15_468 ();
 sg13g2_decap_4 FILLER_15_475 ();
 sg13g2_fill_1 FILLER_15_485 ();
 sg13g2_decap_4 FILLER_15_500 ();
 sg13g2_fill_2 FILLER_15_504 ();
 sg13g2_fill_2 FILLER_15_578 ();
 sg13g2_fill_1 FILLER_15_580 ();
 sg13g2_fill_2 FILLER_15_613 ();
 sg13g2_decap_4 FILLER_15_635 ();
 sg13g2_fill_1 FILLER_15_639 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_fill_2 FILLER_15_669 ();
 sg13g2_fill_1 FILLER_15_671 ();
 sg13g2_fill_2 FILLER_15_708 ();
 sg13g2_fill_1 FILLER_15_710 ();
 sg13g2_fill_2 FILLER_15_720 ();
 sg13g2_decap_4 FILLER_15_727 ();
 sg13g2_fill_2 FILLER_15_731 ();
 sg13g2_fill_1 FILLER_15_741 ();
 sg13g2_decap_4 FILLER_15_755 ();
 sg13g2_fill_1 FILLER_15_759 ();
 sg13g2_fill_1 FILLER_15_794 ();
 sg13g2_fill_1 FILLER_15_799 ();
 sg13g2_fill_2 FILLER_15_814 ();
 sg13g2_decap_8 FILLER_15_824 ();
 sg13g2_fill_2 FILLER_15_831 ();
 sg13g2_fill_2 FILLER_15_842 ();
 sg13g2_fill_2 FILLER_15_856 ();
 sg13g2_fill_2 FILLER_15_863 ();
 sg13g2_fill_1 FILLER_15_893 ();
 sg13g2_fill_2 FILLER_15_969 ();
 sg13g2_fill_2 FILLER_15_1027 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_38 ();
 sg13g2_fill_2 FILLER_16_45 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_decap_4 FILLER_16_190 ();
 sg13g2_decap_8 FILLER_16_215 ();
 sg13g2_decap_8 FILLER_16_222 ();
 sg13g2_decap_4 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_260 ();
 sg13g2_decap_4 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_fill_2 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_315 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_379 ();
 sg13g2_fill_2 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_1 FILLER_16_430 ();
 sg13g2_fill_2 FILLER_16_440 ();
 sg13g2_fill_1 FILLER_16_473 ();
 sg13g2_decap_8 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_521 ();
 sg13g2_decap_4 FILLER_16_528 ();
 sg13g2_decap_8 FILLER_16_541 ();
 sg13g2_fill_2 FILLER_16_548 ();
 sg13g2_fill_1 FILLER_16_550 ();
 sg13g2_fill_1 FILLER_16_565 ();
 sg13g2_fill_1 FILLER_16_580 ();
 sg13g2_decap_4 FILLER_16_589 ();
 sg13g2_decap_8 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_604 ();
 sg13g2_fill_1 FILLER_16_619 ();
 sg13g2_decap_4 FILLER_16_628 ();
 sg13g2_fill_1 FILLER_16_632 ();
 sg13g2_fill_2 FILLER_16_675 ();
 sg13g2_fill_2 FILLER_16_690 ();
 sg13g2_fill_1 FILLER_16_692 ();
 sg13g2_decap_8 FILLER_16_720 ();
 sg13g2_decap_4 FILLER_16_727 ();
 sg13g2_fill_1 FILLER_16_731 ();
 sg13g2_decap_8 FILLER_16_744 ();
 sg13g2_decap_8 FILLER_16_751 ();
 sg13g2_decap_8 FILLER_16_758 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_fill_1 FILLER_16_767 ();
 sg13g2_fill_1 FILLER_16_772 ();
 sg13g2_decap_4 FILLER_16_779 ();
 sg13g2_fill_2 FILLER_16_807 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_fill_2 FILLER_16_837 ();
 sg13g2_fill_1 FILLER_16_839 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_fill_2 FILLER_16_851 ();
 sg13g2_fill_1 FILLER_16_853 ();
 sg13g2_fill_1 FILLER_16_859 ();
 sg13g2_fill_2 FILLER_16_892 ();
 sg13g2_fill_1 FILLER_16_894 ();
 sg13g2_decap_8 FILLER_16_904 ();
 sg13g2_decap_4 FILLER_16_911 ();
 sg13g2_decap_8 FILLER_16_936 ();
 sg13g2_decap_8 FILLER_16_943 ();
 sg13g2_decap_8 FILLER_16_950 ();
 sg13g2_decap_8 FILLER_16_957 ();
 sg13g2_decap_8 FILLER_16_964 ();
 sg13g2_decap_4 FILLER_16_971 ();
 sg13g2_fill_2 FILLER_16_992 ();
 sg13g2_decap_8 FILLER_16_1020 ();
 sg13g2_fill_2 FILLER_16_1027 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_decap_4 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_fill_1 FILLER_17_247 ();
 sg13g2_decap_4 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_271 ();
 sg13g2_decap_8 FILLER_17_285 ();
 sg13g2_fill_2 FILLER_17_292 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_decap_4 FILLER_17_299 ();
 sg13g2_fill_2 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_fill_1 FILLER_17_407 ();
 sg13g2_fill_2 FILLER_17_435 ();
 sg13g2_fill_1 FILLER_17_437 ();
 sg13g2_fill_1 FILLER_17_442 ();
 sg13g2_fill_2 FILLER_17_447 ();
 sg13g2_fill_2 FILLER_17_455 ();
 sg13g2_fill_2 FILLER_17_470 ();
 sg13g2_fill_1 FILLER_17_505 ();
 sg13g2_fill_1 FILLER_17_537 ();
 sg13g2_fill_2 FILLER_17_551 ();
 sg13g2_decap_8 FILLER_17_580 ();
 sg13g2_fill_1 FILLER_17_587 ();
 sg13g2_decap_8 FILLER_17_625 ();
 sg13g2_decap_8 FILLER_17_632 ();
 sg13g2_fill_2 FILLER_17_639 ();
 sg13g2_fill_2 FILLER_17_645 ();
 sg13g2_fill_1 FILLER_17_666 ();
 sg13g2_fill_1 FILLER_17_680 ();
 sg13g2_fill_2 FILLER_17_694 ();
 sg13g2_fill_2 FILLER_17_700 ();
 sg13g2_fill_1 FILLER_17_702 ();
 sg13g2_decap_8 FILLER_17_716 ();
 sg13g2_decap_4 FILLER_17_723 ();
 sg13g2_fill_2 FILLER_17_737 ();
 sg13g2_fill_1 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_fill_1 FILLER_17_784 ();
 sg13g2_fill_2 FILLER_17_790 ();
 sg13g2_fill_1 FILLER_17_800 ();
 sg13g2_fill_2 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_827 ();
 sg13g2_decap_8 FILLER_17_834 ();
 sg13g2_decap_8 FILLER_17_841 ();
 sg13g2_fill_2 FILLER_17_848 ();
 sg13g2_fill_1 FILLER_17_850 ();
 sg13g2_fill_2 FILLER_17_857 ();
 sg13g2_fill_1 FILLER_17_859 ();
 sg13g2_fill_2 FILLER_17_877 ();
 sg13g2_decap_8 FILLER_17_900 ();
 sg13g2_decap_8 FILLER_17_907 ();
 sg13g2_decap_4 FILLER_17_914 ();
 sg13g2_decap_8 FILLER_17_933 ();
 sg13g2_decap_8 FILLER_17_940 ();
 sg13g2_decap_4 FILLER_17_965 ();
 sg13g2_fill_2 FILLER_17_969 ();
 sg13g2_fill_1 FILLER_17_1000 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_fill_1 FILLER_18_27 ();
 sg13g2_decap_8 FILLER_18_33 ();
 sg13g2_fill_2 FILLER_18_40 ();
 sg13g2_decap_4 FILLER_18_46 ();
 sg13g2_fill_2 FILLER_18_90 ();
 sg13g2_fill_1 FILLER_18_92 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_2 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_141 ();
 sg13g2_decap_4 FILLER_18_197 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_fill_1 FILLER_18_254 ();
 sg13g2_fill_2 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_4 FILLER_18_300 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_fill_2 FILLER_18_330 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_fill_2 FILLER_18_383 ();
 sg13g2_decap_4 FILLER_18_427 ();
 sg13g2_fill_2 FILLER_18_435 ();
 sg13g2_decap_4 FILLER_18_443 ();
 sg13g2_fill_2 FILLER_18_447 ();
 sg13g2_fill_1 FILLER_18_462 ();
 sg13g2_fill_1 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_4 FILLER_18_521 ();
 sg13g2_fill_2 FILLER_18_525 ();
 sg13g2_fill_2 FILLER_18_562 ();
 sg13g2_decap_8 FILLER_18_596 ();
 sg13g2_fill_2 FILLER_18_603 ();
 sg13g2_decap_8 FILLER_18_622 ();
 sg13g2_decap_4 FILLER_18_629 ();
 sg13g2_fill_2 FILLER_18_633 ();
 sg13g2_fill_2 FILLER_18_650 ();
 sg13g2_decap_4 FILLER_18_675 ();
 sg13g2_fill_2 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_fill_2 FILLER_18_728 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_fill_2 FILLER_18_760 ();
 sg13g2_decap_4 FILLER_18_789 ();
 sg13g2_fill_1 FILLER_18_793 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_fill_2 FILLER_18_852 ();
 sg13g2_fill_1 FILLER_18_854 ();
 sg13g2_fill_2 FILLER_18_902 ();
 sg13g2_fill_1 FILLER_18_904 ();
 sg13g2_fill_2 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_1020 ();
 sg13g2_fill_2 FILLER_18_1027 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_15 ();
 sg13g2_fill_1 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_decap_4 FILLER_19_41 ();
 sg13g2_decap_4 FILLER_19_50 ();
 sg13g2_decap_4 FILLER_19_67 ();
 sg13g2_fill_2 FILLER_19_71 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_decap_4 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_173 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_2 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_4 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_356 ();
 sg13g2_decap_4 FILLER_19_363 ();
 sg13g2_decap_4 FILLER_19_373 ();
 sg13g2_fill_2 FILLER_19_377 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_fill_1 FILLER_19_404 ();
 sg13g2_decap_8 FILLER_19_409 ();
 sg13g2_decap_4 FILLER_19_416 ();
 sg13g2_fill_2 FILLER_19_420 ();
 sg13g2_fill_1 FILLER_19_435 ();
 sg13g2_fill_2 FILLER_19_467 ();
 sg13g2_fill_1 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_487 ();
 sg13g2_decap_8 FILLER_19_494 ();
 sg13g2_fill_1 FILLER_19_501 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_fill_1 FILLER_19_531 ();
 sg13g2_decap_4 FILLER_19_545 ();
 sg13g2_fill_1 FILLER_19_549 ();
 sg13g2_fill_1 FILLER_19_580 ();
 sg13g2_fill_2 FILLER_19_616 ();
 sg13g2_fill_2 FILLER_19_645 ();
 sg13g2_fill_1 FILLER_19_647 ();
 sg13g2_fill_2 FILLER_19_667 ();
 sg13g2_fill_1 FILLER_19_669 ();
 sg13g2_fill_2 FILLER_19_697 ();
 sg13g2_fill_1 FILLER_19_699 ();
 sg13g2_fill_2 FILLER_19_706 ();
 sg13g2_decap_4 FILLER_19_712 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_fill_2 FILLER_19_732 ();
 sg13g2_fill_1 FILLER_19_734 ();
 sg13g2_decap_4 FILLER_19_744 ();
 sg13g2_fill_2 FILLER_19_780 ();
 sg13g2_fill_1 FILLER_19_782 ();
 sg13g2_decap_4 FILLER_19_792 ();
 sg13g2_fill_2 FILLER_19_809 ();
 sg13g2_fill_2 FILLER_19_834 ();
 sg13g2_fill_1 FILLER_19_836 ();
 sg13g2_decap_4 FILLER_19_846 ();
 sg13g2_fill_1 FILLER_19_858 ();
 sg13g2_decap_4 FILLER_19_871 ();
 sg13g2_fill_1 FILLER_19_893 ();
 sg13g2_fill_2 FILLER_19_919 ();
 sg13g2_fill_1 FILLER_19_921 ();
 sg13g2_decap_8 FILLER_19_938 ();
 sg13g2_fill_2 FILLER_19_945 ();
 sg13g2_fill_1 FILLER_19_947 ();
 sg13g2_fill_2 FILLER_19_966 ();
 sg13g2_fill_2 FILLER_19_978 ();
 sg13g2_fill_1 FILLER_19_980 ();
 sg13g2_fill_2 FILLER_19_1026 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_51 ();
 sg13g2_fill_2 FILLER_20_72 ();
 sg13g2_fill_2 FILLER_20_148 ();
 sg13g2_fill_2 FILLER_20_176 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_decap_4 FILLER_20_281 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_4 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_432 ();
 sg13g2_decap_8 FILLER_20_439 ();
 sg13g2_fill_2 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_462 ();
 sg13g2_fill_2 FILLER_20_473 ();
 sg13g2_decap_4 FILLER_20_518 ();
 sg13g2_decap_4 FILLER_20_527 ();
 sg13g2_fill_2 FILLER_20_531 ();
 sg13g2_fill_2 FILLER_20_551 ();
 sg13g2_fill_1 FILLER_20_553 ();
 sg13g2_decap_4 FILLER_20_567 ();
 sg13g2_fill_1 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_598 ();
 sg13g2_fill_2 FILLER_20_605 ();
 sg13g2_fill_1 FILLER_20_607 ();
 sg13g2_fill_1 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_671 ();
 sg13g2_decap_4 FILLER_20_678 ();
 sg13g2_fill_1 FILLER_20_682 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_fill_2 FILLER_20_728 ();
 sg13g2_fill_1 FILLER_20_730 ();
 sg13g2_fill_2 FILLER_20_735 ();
 sg13g2_fill_1 FILLER_20_745 ();
 sg13g2_fill_1 FILLER_20_752 ();
 sg13g2_fill_1 FILLER_20_784 ();
 sg13g2_fill_2 FILLER_20_804 ();
 sg13g2_fill_1 FILLER_20_806 ();
 sg13g2_fill_2 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_871 ();
 sg13g2_decap_8 FILLER_20_878 ();
 sg13g2_fill_2 FILLER_20_885 ();
 sg13g2_fill_2 FILLER_20_937 ();
 sg13g2_fill_1 FILLER_20_939 ();
 sg13g2_decap_4 FILLER_20_949 ();
 sg13g2_decap_4 FILLER_20_962 ();
 sg13g2_fill_1 FILLER_20_966 ();
 sg13g2_decap_4 FILLER_20_975 ();
 sg13g2_fill_1 FILLER_20_983 ();
 sg13g2_fill_1 FILLER_20_990 ();
 sg13g2_decap_8 FILLER_20_1018 ();
 sg13g2_decap_4 FILLER_20_1025 ();
 sg13g2_fill_2 FILLER_21_27 ();
 sg13g2_fill_2 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_126 ();
 sg13g2_decap_4 FILLER_21_165 ();
 sg13g2_fill_1 FILLER_21_169 ();
 sg13g2_decap_4 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_205 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_2 FILLER_21_218 ();
 sg13g2_decap_4 FILLER_21_264 ();
 sg13g2_fill_2 FILLER_21_299 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_4 FILLER_21_338 ();
 sg13g2_fill_1 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_400 ();
 sg13g2_fill_1 FILLER_21_409 ();
 sg13g2_decap_8 FILLER_21_437 ();
 sg13g2_fill_2 FILLER_21_444 ();
 sg13g2_fill_1 FILLER_21_446 ();
 sg13g2_fill_1 FILLER_21_517 ();
 sg13g2_decap_4 FILLER_21_572 ();
 sg13g2_fill_2 FILLER_21_576 ();
 sg13g2_fill_2 FILLER_21_604 ();
 sg13g2_fill_1 FILLER_21_606 ();
 sg13g2_fill_2 FILLER_21_620 ();
 sg13g2_fill_1 FILLER_21_622 ();
 sg13g2_fill_1 FILLER_21_650 ();
 sg13g2_fill_1 FILLER_21_655 ();
 sg13g2_fill_1 FILLER_21_666 ();
 sg13g2_decap_4 FILLER_21_771 ();
 sg13g2_fill_1 FILLER_21_775 ();
 sg13g2_decap_4 FILLER_21_785 ();
 sg13g2_decap_8 FILLER_21_822 ();
 sg13g2_decap_8 FILLER_21_829 ();
 sg13g2_fill_1 FILLER_21_836 ();
 sg13g2_fill_2 FILLER_21_850 ();
 sg13g2_fill_2 FILLER_21_858 ();
 sg13g2_decap_4 FILLER_21_905 ();
 sg13g2_fill_1 FILLER_21_909 ();
 sg13g2_decap_8 FILLER_21_913 ();
 sg13g2_decap_4 FILLER_21_920 ();
 sg13g2_fill_2 FILLER_21_924 ();
 sg13g2_fill_1 FILLER_21_983 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_4 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_8 ();
 sg13g2_decap_4 FILLER_22_22 ();
 sg13g2_fill_2 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_37 ();
 sg13g2_fill_2 FILLER_22_57 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_142 ();
 sg13g2_decap_8 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_8 FILLER_22_206 ();
 sg13g2_fill_2 FILLER_22_213 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_fill_2 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_281 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_fill_1 FILLER_22_367 ();
 sg13g2_fill_1 FILLER_22_373 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_22_391 ();
 sg13g2_fill_2 FILLER_22_433 ();
 sg13g2_fill_1 FILLER_22_479 ();
 sg13g2_fill_2 FILLER_22_493 ();
 sg13g2_fill_1 FILLER_22_495 ();
 sg13g2_fill_2 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_507 ();
 sg13g2_fill_2 FILLER_22_534 ();
 sg13g2_fill_1 FILLER_22_618 ();
 sg13g2_fill_2 FILLER_22_684 ();
 sg13g2_fill_1 FILLER_22_686 ();
 sg13g2_fill_1 FILLER_22_696 ();
 sg13g2_decap_8 FILLER_22_719 ();
 sg13g2_fill_2 FILLER_22_726 ();
 sg13g2_fill_1 FILLER_22_728 ();
 sg13g2_fill_1 FILLER_22_748 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_4 FILLER_22_781 ();
 sg13g2_fill_1 FILLER_22_785 ();
 sg13g2_fill_1 FILLER_22_807 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_4 FILLER_22_819 ();
 sg13g2_fill_2 FILLER_22_849 ();
 sg13g2_fill_2 FILLER_22_874 ();
 sg13g2_fill_1 FILLER_22_876 ();
 sg13g2_fill_1 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_908 ();
 sg13g2_fill_2 FILLER_22_915 ();
 sg13g2_fill_1 FILLER_22_917 ();
 sg13g2_decap_8 FILLER_22_945 ();
 sg13g2_decap_8 FILLER_22_952 ();
 sg13g2_decap_4 FILLER_22_959 ();
 sg13g2_fill_1 FILLER_22_963 ();
 sg13g2_fill_2 FILLER_22_970 ();
 sg13g2_fill_1 FILLER_22_972 ();
 sg13g2_fill_1 FILLER_22_979 ();
 sg13g2_fill_1 FILLER_22_1001 ();
 sg13g2_fill_2 FILLER_23_33 ();
 sg13g2_decap_8 FILLER_23_48 ();
 sg13g2_decap_4 FILLER_23_55 ();
 sg13g2_decap_4 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_decap_4 FILLER_23_148 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_fill_1 FILLER_23_217 ();
 sg13g2_fill_1 FILLER_23_223 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_4 FILLER_23_302 ();
 sg13g2_fill_2 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_349 ();
 sg13g2_decap_4 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_fill_1 FILLER_23_395 ();
 sg13g2_fill_2 FILLER_23_401 ();
 sg13g2_fill_2 FILLER_23_417 ();
 sg13g2_fill_1 FILLER_23_419 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_fill_2 FILLER_23_465 ();
 sg13g2_fill_1 FILLER_23_467 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_fill_1 FILLER_23_480 ();
 sg13g2_fill_1 FILLER_23_508 ();
 sg13g2_fill_1 FILLER_23_529 ();
 sg13g2_decap_4 FILLER_23_573 ();
 sg13g2_fill_2 FILLER_23_577 ();
 sg13g2_fill_2 FILLER_23_610 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_4 FILLER_23_630 ();
 sg13g2_fill_2 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_659 ();
 sg13g2_fill_2 FILLER_23_666 ();
 sg13g2_fill_1 FILLER_23_668 ();
 sg13g2_fill_2 FILLER_23_682 ();
 sg13g2_fill_1 FILLER_23_688 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_fill_1 FILLER_23_706 ();
 sg13g2_decap_8 FILLER_23_724 ();
 sg13g2_fill_1 FILLER_23_735 ();
 sg13g2_fill_2 FILLER_23_742 ();
 sg13g2_fill_1 FILLER_23_744 ();
 sg13g2_fill_1 FILLER_23_749 ();
 sg13g2_fill_2 FILLER_23_759 ();
 sg13g2_decap_4 FILLER_23_788 ();
 sg13g2_fill_2 FILLER_23_792 ();
 sg13g2_fill_2 FILLER_23_807 ();
 sg13g2_fill_1 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_836 ();
 sg13g2_decap_8 FILLER_23_843 ();
 sg13g2_decap_4 FILLER_23_850 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_fill_2 FILLER_23_896 ();
 sg13g2_fill_1 FILLER_23_898 ();
 sg13g2_fill_1 FILLER_23_940 ();
 sg13g2_decap_8 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_952 ();
 sg13g2_decap_4 FILLER_23_959 ();
 sg13g2_fill_1 FILLER_23_984 ();
 sg13g2_fill_2 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1018 ();
 sg13g2_decap_4 FILLER_23_1025 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_18 ();
 sg13g2_fill_2 FILLER_24_68 ();
 sg13g2_fill_1 FILLER_24_97 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_113 ();
 sg13g2_fill_1 FILLER_24_117 ();
 sg13g2_decap_4 FILLER_24_121 ();
 sg13g2_decap_4 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_1 FILLER_24_249 ();
 sg13g2_fill_2 FILLER_24_291 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_fill_1 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_4 FILLER_24_431 ();
 sg13g2_fill_2 FILLER_24_435 ();
 sg13g2_decap_4 FILLER_24_450 ();
 sg13g2_fill_1 FILLER_24_454 ();
 sg13g2_decap_4 FILLER_24_480 ();
 sg13g2_fill_1 FILLER_24_484 ();
 sg13g2_fill_1 FILLER_24_502 ();
 sg13g2_decap_4 FILLER_24_530 ();
 sg13g2_fill_2 FILLER_24_534 ();
 sg13g2_fill_2 FILLER_24_555 ();
 sg13g2_fill_1 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_fill_2 FILLER_24_571 ();
 sg13g2_fill_1 FILLER_24_573 ();
 sg13g2_fill_2 FILLER_24_584 ();
 sg13g2_decap_4 FILLER_24_644 ();
 sg13g2_fill_1 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_668 ();
 sg13g2_decap_4 FILLER_24_675 ();
 sg13g2_fill_1 FILLER_24_687 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_fill_2 FILLER_24_788 ();
 sg13g2_fill_1 FILLER_24_790 ();
 sg13g2_fill_1 FILLER_24_804 ();
 sg13g2_decap_8 FILLER_24_818 ();
 sg13g2_decap_4 FILLER_24_825 ();
 sg13g2_fill_2 FILLER_24_829 ();
 sg13g2_fill_1 FILLER_24_844 ();
 sg13g2_fill_1 FILLER_24_861 ();
 sg13g2_decap_8 FILLER_24_888 ();
 sg13g2_fill_2 FILLER_24_895 ();
 sg13g2_decap_4 FILLER_24_935 ();
 sg13g2_fill_1 FILLER_24_939 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_fill_2 FILLER_25_69 ();
 sg13g2_fill_2 FILLER_25_90 ();
 sg13g2_fill_1 FILLER_25_92 ();
 sg13g2_decap_4 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_106 ();
 sg13g2_decap_8 FILLER_25_122 ();
 sg13g2_decap_8 FILLER_25_129 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_8 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_157 ();
 sg13g2_decap_4 FILLER_25_173 ();
 sg13g2_decap_4 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_261 ();
 sg13g2_decap_8 FILLER_25_292 ();
 sg13g2_fill_1 FILLER_25_348 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_fill_2 FILLER_25_426 ();
 sg13g2_fill_1 FILLER_25_428 ();
 sg13g2_fill_2 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_523 ();
 sg13g2_fill_2 FILLER_25_530 ();
 sg13g2_fill_2 FILLER_25_537 ();
 sg13g2_fill_1 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_555 ();
 sg13g2_decap_8 FILLER_25_562 ();
 sg13g2_fill_2 FILLER_25_569 ();
 sg13g2_decap_8 FILLER_25_617 ();
 sg13g2_decap_4 FILLER_25_624 ();
 sg13g2_fill_1 FILLER_25_628 ();
 sg13g2_decap_4 FILLER_25_634 ();
 sg13g2_fill_2 FILLER_25_638 ();
 sg13g2_fill_1 FILLER_25_645 ();
 sg13g2_fill_1 FILLER_25_683 ();
 sg13g2_decap_4 FILLER_25_692 ();
 sg13g2_fill_1 FILLER_25_696 ();
 sg13g2_decap_8 FILLER_25_724 ();
 sg13g2_fill_2 FILLER_25_731 ();
 sg13g2_decap_4 FILLER_25_743 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_785 ();
 sg13g2_fill_2 FILLER_25_792 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_fill_2 FILLER_25_821 ();
 sg13g2_fill_1 FILLER_25_823 ();
 sg13g2_fill_1 FILLER_25_861 ();
 sg13g2_decap_4 FILLER_25_889 ();
 sg13g2_fill_1 FILLER_25_897 ();
 sg13g2_fill_2 FILLER_25_930 ();
 sg13g2_fill_1 FILLER_25_932 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_4 FILLER_25_973 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_48 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_1 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_4 FILLER_26_207 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_292 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_310 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_decap_4 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_decap_4 FILLER_26_376 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_decap_4 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_4 FILLER_26_431 ();
 sg13g2_decap_8 FILLER_26_449 ();
 sg13g2_decap_4 FILLER_26_470 ();
 sg13g2_fill_1 FILLER_26_501 ();
 sg13g2_decap_8 FILLER_26_515 ();
 sg13g2_fill_1 FILLER_26_536 ();
 sg13g2_fill_2 FILLER_26_561 ();
 sg13g2_fill_2 FILLER_26_579 ();
 sg13g2_fill_1 FILLER_26_612 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_4 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_4 FILLER_26_729 ();
 sg13g2_decap_4 FILLER_26_752 ();
 sg13g2_fill_2 FILLER_26_783 ();
 sg13g2_fill_1 FILLER_26_785 ();
 sg13g2_fill_2 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_815 ();
 sg13g2_decap_8 FILLER_26_822 ();
 sg13g2_fill_2 FILLER_26_829 ();
 sg13g2_fill_1 FILLER_26_831 ();
 sg13g2_fill_1 FILLER_26_836 ();
 sg13g2_decap_8 FILLER_26_963 ();
 sg13g2_decap_8 FILLER_26_970 ();
 sg13g2_fill_1 FILLER_26_987 ();
 sg13g2_fill_1 FILLER_26_996 ();
 sg13g2_decap_8 FILLER_26_1019 ();
 sg13g2_fill_2 FILLER_26_1026 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_79 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_4 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_fill_1 FILLER_27_172 ();
 sg13g2_fill_2 FILLER_27_227 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_292 ();
 sg13g2_decap_8 FILLER_27_299 ();
 sg13g2_decap_4 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_310 ();
 sg13g2_decap_4 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_357 ();
 sg13g2_decap_4 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_366 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_435 ();
 sg13g2_fill_1 FILLER_27_437 ();
 sg13g2_decap_8 FILLER_27_451 ();
 sg13g2_fill_2 FILLER_27_458 ();
 sg13g2_fill_1 FILLER_27_460 ();
 sg13g2_decap_4 FILLER_27_491 ();
 sg13g2_fill_1 FILLER_27_495 ();
 sg13g2_fill_1 FILLER_27_523 ();
 sg13g2_fill_2 FILLER_27_533 ();
 sg13g2_fill_1 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_593 ();
 sg13g2_fill_1 FILLER_27_598 ();
 sg13g2_fill_2 FILLER_27_626 ();
 sg13g2_fill_1 FILLER_27_628 ();
 sg13g2_fill_2 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_689 ();
 sg13g2_fill_2 FILLER_27_696 ();
 sg13g2_fill_1 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_4 FILLER_27_723 ();
 sg13g2_fill_2 FILLER_27_727 ();
 sg13g2_fill_1 FILLER_27_756 ();
 sg13g2_fill_2 FILLER_27_781 ();
 sg13g2_fill_1 FILLER_27_866 ();
 sg13g2_fill_1 FILLER_27_875 ();
 sg13g2_fill_1 FILLER_27_888 ();
 sg13g2_decap_8 FILLER_27_900 ();
 sg13g2_decap_4 FILLER_27_907 ();
 sg13g2_fill_2 FILLER_27_911 ();
 sg13g2_fill_2 FILLER_27_988 ();
 sg13g2_fill_2 FILLER_27_1026 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_100 ();
 sg13g2_fill_2 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_246 ();
 sg13g2_fill_2 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_351 ();
 sg13g2_fill_2 FILLER_28_396 ();
 sg13g2_decap_8 FILLER_28_407 ();
 sg13g2_fill_1 FILLER_28_414 ();
 sg13g2_decap_4 FILLER_28_421 ();
 sg13g2_fill_1 FILLER_28_447 ();
 sg13g2_decap_8 FILLER_28_475 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_fill_1 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_fill_2 FILLER_28_553 ();
 sg13g2_fill_2 FILLER_28_581 ();
 sg13g2_fill_2 FILLER_28_610 ();
 sg13g2_fill_2 FILLER_28_652 ();
 sg13g2_fill_1 FILLER_28_694 ();
 sg13g2_decap_4 FILLER_28_726 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_4 FILLER_28_762 ();
 sg13g2_fill_2 FILLER_28_766 ();
 sg13g2_fill_1 FILLER_28_799 ();
 sg13g2_decap_8 FILLER_28_829 ();
 sg13g2_decap_4 FILLER_28_836 ();
 sg13g2_fill_2 FILLER_28_904 ();
 sg13g2_decap_8 FILLER_28_932 ();
 sg13g2_decap_4 FILLER_28_939 ();
 sg13g2_fill_1 FILLER_28_943 ();
 sg13g2_fill_1 FILLER_28_949 ();
 sg13g2_decap_8 FILLER_28_961 ();
 sg13g2_decap_4 FILLER_28_968 ();
 sg13g2_fill_1 FILLER_28_972 ();
 sg13g2_decap_8 FILLER_28_1018 ();
 sg13g2_decap_4 FILLER_28_1025 ();
 sg13g2_decap_4 FILLER_29_4 ();
 sg13g2_fill_1 FILLER_29_8 ();
 sg13g2_fill_1 FILLER_29_38 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_fill_2 FILLER_29_112 ();
 sg13g2_fill_2 FILLER_29_127 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_decap_4 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_232 ();
 sg13g2_decap_8 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_2 FILLER_29_356 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_391 ();
 sg13g2_fill_2 FILLER_29_395 ();
 sg13g2_fill_1 FILLER_29_404 ();
 sg13g2_decap_8 FILLER_29_414 ();
 sg13g2_fill_1 FILLER_29_421 ();
 sg13g2_decap_4 FILLER_29_449 ();
 sg13g2_fill_1 FILLER_29_453 ();
 sg13g2_decap_8 FILLER_29_467 ();
 sg13g2_fill_1 FILLER_29_483 ();
 sg13g2_decap_4 FILLER_29_537 ();
 sg13g2_decap_8 FILLER_29_545 ();
 sg13g2_decap_4 FILLER_29_552 ();
 sg13g2_fill_1 FILLER_29_556 ();
 sg13g2_fill_2 FILLER_29_596 ();
 sg13g2_fill_2 FILLER_29_602 ();
 sg13g2_fill_2 FILLER_29_630 ();
 sg13g2_fill_1 FILLER_29_632 ();
 sg13g2_fill_2 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_fill_2 FILLER_29_729 ();
 sg13g2_fill_1 FILLER_29_731 ();
 sg13g2_decap_8 FILLER_29_745 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_fill_2 FILLER_29_852 ();
 sg13g2_decap_4 FILLER_29_860 ();
 sg13g2_fill_2 FILLER_29_873 ();
 sg13g2_fill_2 FILLER_29_889 ();
 sg13g2_fill_2 FILLER_29_904 ();
 sg13g2_fill_1 FILLER_29_919 ();
 sg13g2_decap_8 FILLER_29_933 ();
 sg13g2_fill_2 FILLER_29_940 ();
 sg13g2_fill_1 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_968 ();
 sg13g2_fill_2 FILLER_29_975 ();
 sg13g2_fill_2 FILLER_29_981 ();
 sg13g2_fill_1 FILLER_29_987 ();
 sg13g2_decap_4 FILLER_29_1024 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_fill_1 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_179 ();
 sg13g2_decap_4 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_243 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_1 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_fill_2 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_4 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_383 ();
 sg13g2_fill_1 FILLER_30_417 ();
 sg13g2_fill_1 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_445 ();
 sg13g2_decap_8 FILLER_30_452 ();
 sg13g2_decap_4 FILLER_30_459 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_4 FILLER_30_497 ();
 sg13g2_fill_1 FILLER_30_501 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_4 FILLER_30_518 ();
 sg13g2_fill_1 FILLER_30_522 ();
 sg13g2_decap_4 FILLER_30_562 ();
 sg13g2_fill_1 FILLER_30_579 ();
 sg13g2_fill_2 FILLER_30_610 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_1 FILLER_30_641 ();
 sg13g2_fill_2 FILLER_30_678 ();
 sg13g2_fill_1 FILLER_30_680 ();
 sg13g2_fill_2 FILLER_30_696 ();
 sg13g2_fill_1 FILLER_30_738 ();
 sg13g2_fill_1 FILLER_30_766 ();
 sg13g2_fill_1 FILLER_30_784 ();
 sg13g2_fill_2 FILLER_30_806 ();
 sg13g2_fill_1 FILLER_30_808 ();
 sg13g2_decap_8 FILLER_30_818 ();
 sg13g2_decap_8 FILLER_30_825 ();
 sg13g2_decap_4 FILLER_30_832 ();
 sg13g2_fill_2 FILLER_30_840 ();
 sg13g2_fill_1 FILLER_30_842 ();
 sg13g2_fill_1 FILLER_30_860 ();
 sg13g2_fill_2 FILLER_30_888 ();
 sg13g2_fill_1 FILLER_30_890 ();
 sg13g2_fill_1 FILLER_30_917 ();
 sg13g2_fill_1 FILLER_30_972 ();
 sg13g2_fill_1 FILLER_30_992 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_68 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_4 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_167 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_decap_4 FILLER_31_215 ();
 sg13g2_decap_4 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_236 ();
 sg13g2_decap_4 FILLER_31_277 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_fill_1 FILLER_31_430 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_503 ();
 sg13g2_fill_1 FILLER_31_510 ();
 sg13g2_decap_8 FILLER_31_545 ();
 sg13g2_decap_8 FILLER_31_552 ();
 sg13g2_fill_2 FILLER_31_559 ();
 sg13g2_fill_1 FILLER_31_561 ();
 sg13g2_decap_4 FILLER_31_598 ();
 sg13g2_fill_1 FILLER_31_615 ();
 sg13g2_fill_2 FILLER_31_722 ();
 sg13g2_fill_1 FILLER_31_724 ();
 sg13g2_fill_1 FILLER_31_792 ();
 sg13g2_fill_2 FILLER_31_822 ();
 sg13g2_fill_1 FILLER_31_824 ();
 sg13g2_fill_1 FILLER_31_842 ();
 sg13g2_fill_2 FILLER_31_888 ();
 sg13g2_fill_2 FILLER_31_895 ();
 sg13g2_fill_1 FILLER_31_897 ();
 sg13g2_decap_4 FILLER_31_929 ();
 sg13g2_fill_2 FILLER_31_933 ();
 sg13g2_decap_8 FILLER_31_948 ();
 sg13g2_decap_8 FILLER_31_955 ();
 sg13g2_decap_8 FILLER_31_962 ();
 sg13g2_fill_1 FILLER_31_969 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_fill_2 FILLER_32_189 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_1 FILLER_32_223 ();
 sg13g2_decap_4 FILLER_32_230 ();
 sg13g2_fill_2 FILLER_32_234 ();
 sg13g2_decap_4 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_301 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_fill_1 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_404 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_fill_2 FILLER_32_490 ();
 sg13g2_fill_1 FILLER_32_519 ();
 sg13g2_fill_1 FILLER_32_528 ();
 sg13g2_decap_8 FILLER_32_556 ();
 sg13g2_decap_4 FILLER_32_563 ();
 sg13g2_fill_1 FILLER_32_567 ();
 sg13g2_decap_4 FILLER_32_608 ();
 sg13g2_fill_2 FILLER_32_659 ();
 sg13g2_fill_1 FILLER_32_661 ();
 sg13g2_decap_4 FILLER_32_668 ();
 sg13g2_fill_1 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_681 ();
 sg13g2_decap_8 FILLER_32_688 ();
 sg13g2_decap_8 FILLER_32_695 ();
 sg13g2_fill_2 FILLER_32_702 ();
 sg13g2_fill_2 FILLER_32_712 ();
 sg13g2_fill_2 FILLER_32_727 ();
 sg13g2_fill_2 FILLER_32_791 ();
 sg13g2_decap_4 FILLER_32_837 ();
 sg13g2_fill_2 FILLER_32_841 ();
 sg13g2_fill_2 FILLER_32_849 ();
 sg13g2_fill_1 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_856 ();
 sg13g2_decap_4 FILLER_32_863 ();
 sg13g2_decap_4 FILLER_32_876 ();
 sg13g2_decap_4 FILLER_32_889 ();
 sg13g2_fill_1 FILLER_32_909 ();
 sg13g2_decap_8 FILLER_32_928 ();
 sg13g2_fill_1 FILLER_32_935 ();
 sg13g2_fill_2 FILLER_32_945 ();
 sg13g2_fill_1 FILLER_32_947 ();
 sg13g2_decap_8 FILLER_32_965 ();
 sg13g2_decap_4 FILLER_32_994 ();
 sg13g2_decap_4 FILLER_32_1025 ();
 sg13g2_fill_2 FILLER_33_27 ();
 sg13g2_fill_2 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_51 ();
 sg13g2_fill_1 FILLER_33_116 ();
 sg13g2_fill_2 FILLER_33_179 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_decap_4 FILLER_33_237 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_1 FILLER_33_269 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_371 ();
 sg13g2_fill_1 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_decap_4 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_33_411 ();
 sg13g2_fill_2 FILLER_33_425 ();
 sg13g2_fill_1 FILLER_33_427 ();
 sg13g2_fill_2 FILLER_33_441 ();
 sg13g2_fill_2 FILLER_33_456 ();
 sg13g2_fill_1 FILLER_33_458 ();
 sg13g2_decap_8 FILLER_33_486 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_fill_2 FILLER_33_507 ();
 sg13g2_fill_1 FILLER_33_509 ();
 sg13g2_fill_2 FILLER_33_519 ();
 sg13g2_fill_1 FILLER_33_521 ();
 sg13g2_decap_8 FILLER_33_531 ();
 sg13g2_decap_8 FILLER_33_538 ();
 sg13g2_decap_8 FILLER_33_545 ();
 sg13g2_fill_2 FILLER_33_552 ();
 sg13g2_fill_1 FILLER_33_554 ();
 sg13g2_decap_8 FILLER_33_610 ();
 sg13g2_fill_2 FILLER_33_677 ();
 sg13g2_fill_1 FILLER_33_679 ();
 sg13g2_decap_4 FILLER_33_686 ();
 sg13g2_fill_2 FILLER_33_690 ();
 sg13g2_decap_4 FILLER_33_718 ();
 sg13g2_fill_2 FILLER_33_722 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_fill_1 FILLER_33_755 ();
 sg13g2_fill_1 FILLER_33_791 ();
 sg13g2_decap_4 FILLER_33_830 ();
 sg13g2_decap_8 FILLER_33_838 ();
 sg13g2_decap_8 FILLER_33_845 ();
 sg13g2_decap_8 FILLER_33_852 ();
 sg13g2_decap_4 FILLER_33_859 ();
 sg13g2_fill_1 FILLER_33_884 ();
 sg13g2_fill_1 FILLER_33_898 ();
 sg13g2_decap_8 FILLER_33_939 ();
 sg13g2_fill_2 FILLER_33_960 ();
 sg13g2_decap_8 FILLER_33_1014 ();
 sg13g2_decap_8 FILLER_33_1021 ();
 sg13g2_fill_1 FILLER_33_1028 ();
 sg13g2_fill_1 FILLER_34_42 ();
 sg13g2_decap_4 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_decap_8 FILLER_34_64 ();
 sg13g2_fill_2 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_decap_4 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_252 ();
 sg13g2_fill_2 FILLER_34_280 ();
 sg13g2_decap_4 FILLER_34_309 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_2 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_426 ();
 sg13g2_fill_2 FILLER_34_463 ();
 sg13g2_decap_4 FILLER_34_492 ();
 sg13g2_fill_1 FILLER_34_496 ();
 sg13g2_fill_2 FILLER_34_510 ();
 sg13g2_fill_1 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_fill_1 FILLER_34_546 ();
 sg13g2_decap_4 FILLER_34_571 ();
 sg13g2_fill_2 FILLER_34_575 ();
 sg13g2_decap_4 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_720 ();
 sg13g2_fill_2 FILLER_34_727 ();
 sg13g2_fill_2 FILLER_34_760 ();
 sg13g2_fill_2 FILLER_34_799 ();
 sg13g2_fill_1 FILLER_34_828 ();
 sg13g2_fill_1 FILLER_34_833 ();
 sg13g2_fill_1 FILLER_34_870 ();
 sg13g2_decap_4 FILLER_34_904 ();
 sg13g2_fill_1 FILLER_34_908 ();
 sg13g2_decap_8 FILLER_34_933 ();
 sg13g2_fill_1 FILLER_34_940 ();
 sg13g2_fill_1 FILLER_34_974 ();
 sg13g2_decap_4 FILLER_34_992 ();
 sg13g2_fill_2 FILLER_34_996 ();
 sg13g2_decap_8 FILLER_34_1007 ();
 sg13g2_decap_8 FILLER_34_1014 ();
 sg13g2_decap_8 FILLER_34_1021 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_35_8 ();
 sg13g2_fill_1 FILLER_35_15 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_1 FILLER_35_81 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_decap_4 FILLER_35_132 ();
 sg13g2_fill_1 FILLER_35_136 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_356 ();
 sg13g2_decap_4 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_471 ();
 sg13g2_fill_2 FILLER_35_498 ();
 sg13g2_fill_1 FILLER_35_500 ();
 sg13g2_fill_1 FILLER_35_528 ();
 sg13g2_decap_8 FILLER_35_572 ();
 sg13g2_decap_4 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_656 ();
 sg13g2_fill_1 FILLER_35_658 ();
 sg13g2_fill_1 FILLER_35_680 ();
 sg13g2_decap_4 FILLER_35_694 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_fill_2 FILLER_35_768 ();
 sg13g2_fill_2 FILLER_35_775 ();
 sg13g2_fill_1 FILLER_35_777 ();
 sg13g2_fill_2 FILLER_35_812 ();
 sg13g2_fill_1 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_829 ();
 sg13g2_decap_4 FILLER_35_836 ();
 sg13g2_fill_1 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_886 ();
 sg13g2_decap_4 FILLER_35_893 ();
 sg13g2_fill_2 FILLER_35_897 ();
 sg13g2_fill_1 FILLER_35_903 ();
 sg13g2_decap_4 FILLER_35_926 ();
 sg13g2_fill_1 FILLER_35_930 ();
 sg13g2_fill_2 FILLER_35_944 ();
 sg13g2_decap_4 FILLER_35_956 ();
 sg13g2_fill_2 FILLER_35_1000 ();
 sg13g2_fill_1 FILLER_35_1002 ();
 sg13g2_decap_8 FILLER_35_1016 ();
 sg13g2_decap_4 FILLER_35_1023 ();
 sg13g2_fill_2 FILLER_35_1027 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_decap_4 FILLER_36_165 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_206 ();
 sg13g2_decap_4 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_237 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_decap_4 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_355 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_394 ();
 sg13g2_fill_2 FILLER_36_408 ();
 sg13g2_fill_2 FILLER_36_423 ();
 sg13g2_fill_1 FILLER_36_425 ();
 sg13g2_decap_4 FILLER_36_438 ();
 sg13g2_decap_4 FILLER_36_465 ();
 sg13g2_fill_1 FILLER_36_469 ();
 sg13g2_decap_4 FILLER_36_478 ();
 sg13g2_fill_1 FILLER_36_482 ();
 sg13g2_decap_4 FILLER_36_488 ();
 sg13g2_decap_4 FILLER_36_498 ();
 sg13g2_fill_2 FILLER_36_519 ();
 sg13g2_fill_1 FILLER_36_521 ();
 sg13g2_fill_2 FILLER_36_544 ();
 sg13g2_fill_1 FILLER_36_546 ();
 sg13g2_fill_1 FILLER_36_559 ();
 sg13g2_decap_8 FILLER_36_569 ();
 sg13g2_fill_1 FILLER_36_589 ();
 sg13g2_decap_4 FILLER_36_598 ();
 sg13g2_fill_1 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_680 ();
 sg13g2_fill_1 FILLER_36_687 ();
 sg13g2_decap_4 FILLER_36_701 ();
 sg13g2_fill_1 FILLER_36_705 ();
 sg13g2_fill_2 FILLER_36_719 ();
 sg13g2_fill_2 FILLER_36_783 ();
 sg13g2_fill_1 FILLER_36_785 ();
 sg13g2_fill_2 FILLER_36_807 ();
 sg13g2_fill_1 FILLER_36_809 ();
 sg13g2_fill_1 FILLER_36_823 ();
 sg13g2_fill_2 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_862 ();
 sg13g2_decap_4 FILLER_36_869 ();
 sg13g2_fill_2 FILLER_36_873 ();
 sg13g2_fill_2 FILLER_36_888 ();
 sg13g2_fill_1 FILLER_36_890 ();
 sg13g2_decap_4 FILLER_36_928 ();
 sg13g2_fill_2 FILLER_36_945 ();
 sg13g2_fill_1 FILLER_36_960 ();
 sg13g2_fill_1 FILLER_36_974 ();
 sg13g2_decap_8 FILLER_36_990 ();
 sg13g2_decap_8 FILLER_36_997 ();
 sg13g2_decap_8 FILLER_36_1004 ();
 sg13g2_decap_8 FILLER_36_1011 ();
 sg13g2_decap_8 FILLER_36_1018 ();
 sg13g2_decap_4 FILLER_36_1025 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_51 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_144 ();
 sg13g2_decap_4 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_328 ();
 sg13g2_fill_2 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_388 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_fill_2 FILLER_37_438 ();
 sg13g2_fill_1 FILLER_37_440 ();
 sg13g2_decap_4 FILLER_37_451 ();
 sg13g2_decap_8 FILLER_37_563 ();
 sg13g2_decap_4 FILLER_37_570 ();
 sg13g2_fill_1 FILLER_37_574 ();
 sg13g2_decap_4 FILLER_37_588 ();
 sg13g2_fill_1 FILLER_37_592 ();
 sg13g2_fill_2 FILLER_37_614 ();
 sg13g2_decap_8 FILLER_37_642 ();
 sg13g2_fill_1 FILLER_37_649 ();
 sg13g2_decap_4 FILLER_37_681 ();
 sg13g2_fill_1 FILLER_37_685 ();
 sg13g2_decap_4 FILLER_37_717 ();
 sg13g2_fill_2 FILLER_37_778 ();
 sg13g2_decap_8 FILLER_37_785 ();
 sg13g2_decap_4 FILLER_37_792 ();
 sg13g2_decap_4 FILLER_37_800 ();
 sg13g2_fill_1 FILLER_37_804 ();
 sg13g2_fill_2 FILLER_37_841 ();
 sg13g2_decap_4 FILLER_37_847 ();
 sg13g2_fill_2 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_885 ();
 sg13g2_decap_4 FILLER_37_892 ();
 sg13g2_fill_1 FILLER_37_896 ();
 sg13g2_fill_2 FILLER_37_926 ();
 sg13g2_fill_1 FILLER_37_928 ();
 sg13g2_fill_2 FILLER_37_968 ();
 sg13g2_decap_8 FILLER_37_1010 ();
 sg13g2_decap_8 FILLER_37_1017 ();
 sg13g2_decap_4 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_30 ();
 sg13g2_fill_1 FILLER_38_50 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_fill_1 FILLER_38_112 ();
 sg13g2_decap_4 FILLER_38_135 ();
 sg13g2_fill_1 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_216 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_246 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_decap_4 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_4 FILLER_38_384 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_fill_1 FILLER_38_434 ();
 sg13g2_decap_4 FILLER_38_452 ();
 sg13g2_fill_2 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_502 ();
 sg13g2_decap_4 FILLER_38_509 ();
 sg13g2_fill_1 FILLER_38_513 ();
 sg13g2_decap_8 FILLER_38_527 ();
 sg13g2_fill_1 FILLER_38_560 ();
 sg13g2_fill_2 FILLER_38_566 ();
 sg13g2_decap_4 FILLER_38_607 ();
 sg13g2_fill_1 FILLER_38_611 ();
 sg13g2_decap_4 FILLER_38_630 ();
 sg13g2_fill_1 FILLER_38_634 ();
 sg13g2_fill_1 FILLER_38_672 ();
 sg13g2_decap_4 FILLER_38_686 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_fill_1 FILLER_38_756 ();
 sg13g2_decap_4 FILLER_38_760 ();
 sg13g2_fill_2 FILLER_38_773 ();
 sg13g2_fill_2 FILLER_38_788 ();
 sg13g2_fill_1 FILLER_38_790 ();
 sg13g2_decap_4 FILLER_38_797 ();
 sg13g2_fill_2 FILLER_38_801 ();
 sg13g2_fill_2 FILLER_38_855 ();
 sg13g2_fill_1 FILLER_38_857 ();
 sg13g2_fill_2 FILLER_38_871 ();
 sg13g2_fill_1 FILLER_38_873 ();
 sg13g2_fill_2 FILLER_38_893 ();
 sg13g2_fill_1 FILLER_38_895 ();
 sg13g2_fill_1 FILLER_38_909 ();
 sg13g2_fill_1 FILLER_38_932 ();
 sg13g2_fill_2 FILLER_38_979 ();
 sg13g2_fill_1 FILLER_38_981 ();
 sg13g2_decap_8 FILLER_38_1009 ();
 sg13g2_decap_8 FILLER_38_1016 ();
 sg13g2_decap_4 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1027 ();
 sg13g2_fill_2 FILLER_39_37 ();
 sg13g2_fill_1 FILLER_39_66 ();
 sg13g2_fill_2 FILLER_39_220 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_fill_1 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_269 ();
 sg13g2_decap_8 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_4 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_332 ();
 sg13g2_fill_1 FILLER_39_334 ();
 sg13g2_fill_2 FILLER_39_352 ();
 sg13g2_fill_1 FILLER_39_354 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_fill_2 FILLER_39_418 ();
 sg13g2_fill_1 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_437 ();
 sg13g2_decap_4 FILLER_39_444 ();
 sg13g2_fill_2 FILLER_39_448 ();
 sg13g2_fill_2 FILLER_39_484 ();
 sg13g2_fill_1 FILLER_39_486 ();
 sg13g2_decap_4 FILLER_39_504 ();
 sg13g2_fill_1 FILLER_39_521 ();
 sg13g2_decap_8 FILLER_39_587 ();
 sg13g2_fill_2 FILLER_39_594 ();
 sg13g2_fill_1 FILLER_39_596 ();
 sg13g2_decap_8 FILLER_39_610 ();
 sg13g2_fill_2 FILLER_39_617 ();
 sg13g2_fill_1 FILLER_39_619 ();
 sg13g2_fill_1 FILLER_39_685 ();
 sg13g2_decap_4 FILLER_39_756 ();
 sg13g2_fill_2 FILLER_39_766 ();
 sg13g2_fill_2 FILLER_39_781 ();
 sg13g2_fill_1 FILLER_39_783 ();
 sg13g2_decap_8 FILLER_39_824 ();
 sg13g2_decap_4 FILLER_39_831 ();
 sg13g2_fill_2 FILLER_39_835 ();
 sg13g2_decap_8 FILLER_39_856 ();
 sg13g2_fill_1 FILLER_39_863 ();
 sg13g2_fill_2 FILLER_39_899 ();
 sg13g2_fill_1 FILLER_39_934 ();
 sg13g2_fill_1 FILLER_39_948 ();
 sg13g2_decap_4 FILLER_39_967 ();
 sg13g2_fill_2 FILLER_39_984 ();
 sg13g2_fill_1 FILLER_39_986 ();
 sg13g2_decap_8 FILLER_39_1005 ();
 sg13g2_decap_8 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1019 ();
 sg13g2_fill_2 FILLER_39_1026 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_1 FILLER_40_30 ();
 sg13g2_fill_1 FILLER_40_37 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_1 FILLER_40_104 ();
 sg13g2_fill_2 FILLER_40_134 ();
 sg13g2_decap_4 FILLER_40_172 ();
 sg13g2_decap_8 FILLER_40_199 ();
 sg13g2_fill_1 FILLER_40_206 ();
 sg13g2_decap_8 FILLER_40_216 ();
 sg13g2_fill_1 FILLER_40_223 ();
 sg13g2_fill_1 FILLER_40_237 ();
 sg13g2_decap_4 FILLER_40_244 ();
 sg13g2_decap_8 FILLER_40_276 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_285 ();
 sg13g2_fill_2 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_fill_2 FILLER_40_331 ();
 sg13g2_fill_1 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_345 ();
 sg13g2_fill_1 FILLER_40_347 ();
 sg13g2_fill_2 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_fill_2 FILLER_40_435 ();
 sg13g2_fill_1 FILLER_40_442 ();
 sg13g2_fill_1 FILLER_40_456 ();
 sg13g2_fill_1 FILLER_40_471 ();
 sg13g2_decap_4 FILLER_40_493 ();
 sg13g2_decap_8 FILLER_40_501 ();
 sg13g2_decap_4 FILLER_40_521 ();
 sg13g2_fill_2 FILLER_40_525 ();
 sg13g2_fill_1 FILLER_40_545 ();
 sg13g2_decap_8 FILLER_40_559 ();
 sg13g2_decap_8 FILLER_40_566 ();
 sg13g2_decap_4 FILLER_40_599 ();
 sg13g2_fill_1 FILLER_40_642 ();
 sg13g2_fill_2 FILLER_40_670 ();
 sg13g2_fill_1 FILLER_40_711 ();
 sg13g2_fill_2 FILLER_40_734 ();
 sg13g2_fill_1 FILLER_40_785 ();
 sg13g2_decap_8 FILLER_40_799 ();
 sg13g2_decap_8 FILLER_40_806 ();
 sg13g2_decap_8 FILLER_40_813 ();
 sg13g2_decap_4 FILLER_40_820 ();
 sg13g2_fill_1 FILLER_40_824 ();
 sg13g2_fill_2 FILLER_40_838 ();
 sg13g2_decap_4 FILLER_40_877 ();
 sg13g2_fill_2 FILLER_40_890 ();
 sg13g2_fill_1 FILLER_40_892 ();
 sg13g2_fill_2 FILLER_40_910 ();
 sg13g2_fill_1 FILLER_40_912 ();
 sg13g2_decap_4 FILLER_40_926 ();
 sg13g2_fill_2 FILLER_40_930 ();
 sg13g2_fill_2 FILLER_40_945 ();
 sg13g2_fill_1 FILLER_40_947 ();
 sg13g2_decap_8 FILLER_40_1019 ();
 sg13g2_fill_2 FILLER_40_1026 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_68 ();
 sg13g2_fill_2 FILLER_41_96 ();
 sg13g2_fill_1 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_131 ();
 sg13g2_decap_4 FILLER_41_170 ();
 sg13g2_fill_2 FILLER_41_174 ();
 sg13g2_decap_4 FILLER_41_189 ();
 sg13g2_fill_2 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_256 ();
 sg13g2_fill_2 FILLER_41_263 ();
 sg13g2_fill_1 FILLER_41_265 ();
 sg13g2_fill_2 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_281 ();
 sg13g2_fill_2 FILLER_41_310 ();
 sg13g2_fill_1 FILLER_41_317 ();
 sg13g2_fill_2 FILLER_41_377 ();
 sg13g2_fill_1 FILLER_41_379 ();
 sg13g2_fill_2 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_432 ();
 sg13g2_fill_1 FILLER_41_461 ();
 sg13g2_fill_1 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_514 ();
 sg13g2_decap_4 FILLER_41_528 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_fill_1 FILLER_41_547 ();
 sg13g2_fill_1 FILLER_41_558 ();
 sg13g2_decap_4 FILLER_41_572 ();
 sg13g2_fill_2 FILLER_41_604 ();
 sg13g2_fill_2 FILLER_41_683 ();
 sg13g2_fill_2 FILLER_41_711 ();
 sg13g2_fill_1 FILLER_41_713 ();
 sg13g2_decap_4 FILLER_41_727 ();
 sg13g2_fill_2 FILLER_41_731 ();
 sg13g2_fill_2 FILLER_41_750 ();
 sg13g2_fill_2 FILLER_41_756 ();
 sg13g2_fill_2 FILLER_41_797 ();
 sg13g2_decap_8 FILLER_41_804 ();
 sg13g2_decap_4 FILLER_41_811 ();
 sg13g2_fill_2 FILLER_41_815 ();
 sg13g2_fill_2 FILLER_41_830 ();
 sg13g2_decap_8 FILLER_41_859 ();
 sg13g2_decap_4 FILLER_41_871 ();
 sg13g2_fill_1 FILLER_41_875 ();
 sg13g2_fill_1 FILLER_41_889 ();
 sg13g2_fill_2 FILLER_41_911 ();
 sg13g2_fill_1 FILLER_41_913 ();
 sg13g2_decap_8 FILLER_41_941 ();
 sg13g2_fill_1 FILLER_41_948 ();
 sg13g2_fill_2 FILLER_41_962 ();
 sg13g2_decap_8 FILLER_41_1018 ();
 sg13g2_decap_4 FILLER_41_1025 ();
 sg13g2_fill_1 FILLER_42_27 ();
 sg13g2_fill_1 FILLER_42_47 ();
 sg13g2_decap_8 FILLER_42_102 ();
 sg13g2_fill_2 FILLER_42_109 ();
 sg13g2_fill_2 FILLER_42_130 ();
 sg13g2_decap_4 FILLER_42_157 ();
 sg13g2_fill_1 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_180 ();
 sg13g2_fill_1 FILLER_42_197 ();
 sg13g2_fill_2 FILLER_42_203 ();
 sg13g2_decap_4 FILLER_42_219 ();
 sg13g2_fill_1 FILLER_42_223 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_249 ();
 sg13g2_decap_8 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_286 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_303 ();
 sg13g2_fill_1 FILLER_42_327 ();
 sg13g2_fill_2 FILLER_42_334 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_decap_4 FILLER_42_354 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_decap_4 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_412 ();
 sg13g2_fill_2 FILLER_42_418 ();
 sg13g2_decap_8 FILLER_42_426 ();
 sg13g2_decap_8 FILLER_42_433 ();
 sg13g2_fill_2 FILLER_42_440 ();
 sg13g2_fill_1 FILLER_42_442 ();
 sg13g2_fill_2 FILLER_42_452 ();
 sg13g2_fill_1 FILLER_42_488 ();
 sg13g2_fill_1 FILLER_42_515 ();
 sg13g2_decap_4 FILLER_42_522 ();
 sg13g2_fill_1 FILLER_42_526 ();
 sg13g2_decap_4 FILLER_42_549 ();
 sg13g2_fill_1 FILLER_42_553 ();
 sg13g2_fill_1 FILLER_42_572 ();
 sg13g2_fill_2 FILLER_42_612 ();
 sg13g2_fill_1 FILLER_42_614 ();
 sg13g2_decap_8 FILLER_42_671 ();
 sg13g2_decap_8 FILLER_42_678 ();
 sg13g2_decap_8 FILLER_42_685 ();
 sg13g2_fill_1 FILLER_42_692 ();
 sg13g2_fill_2 FILLER_42_706 ();
 sg13g2_fill_1 FILLER_42_708 ();
 sg13g2_fill_2 FILLER_42_748 ();
 sg13g2_fill_1 FILLER_42_750 ();
 sg13g2_fill_2 FILLER_42_764 ();
 sg13g2_fill_1 FILLER_42_766 ();
 sg13g2_fill_2 FILLER_42_793 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_decap_8 FILLER_42_840 ();
 sg13g2_fill_1 FILLER_42_847 ();
 sg13g2_fill_2 FILLER_42_872 ();
 sg13g2_fill_2 FILLER_42_887 ();
 sg13g2_fill_1 FILLER_42_889 ();
 sg13g2_decap_4 FILLER_42_911 ();
 sg13g2_fill_1 FILLER_42_929 ();
 sg13g2_fill_2 FILLER_42_957 ();
 sg13g2_fill_1 FILLER_42_959 ();
 sg13g2_decap_4 FILLER_42_964 ();
 sg13g2_fill_1 FILLER_42_968 ();
 sg13g2_fill_1 FILLER_42_985 ();
 sg13g2_decap_8 FILLER_42_1022 ();
 sg13g2_fill_1 FILLER_43_45 ();
 sg13g2_fill_2 FILLER_43_55 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_fill_2 FILLER_43_90 ();
 sg13g2_fill_1 FILLER_43_92 ();
 sg13g2_fill_2 FILLER_43_102 ();
 sg13g2_fill_1 FILLER_43_104 ();
 sg13g2_fill_1 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_164 ();
 sg13g2_decap_8 FILLER_43_183 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_fill_1 FILLER_43_228 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_fill_2 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_279 ();
 sg13g2_fill_2 FILLER_43_317 ();
 sg13g2_fill_1 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_decap_4 FILLER_43_341 ();
 sg13g2_fill_2 FILLER_43_345 ();
 sg13g2_decap_4 FILLER_43_364 ();
 sg13g2_fill_1 FILLER_43_372 ();
 sg13g2_fill_2 FILLER_43_379 ();
 sg13g2_fill_2 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_434 ();
 sg13g2_decap_4 FILLER_43_440 ();
 sg13g2_fill_1 FILLER_43_444 ();
 sg13g2_fill_2 FILLER_43_472 ();
 sg13g2_fill_1 FILLER_43_474 ();
 sg13g2_fill_2 FILLER_43_542 ();
 sg13g2_decap_4 FILLER_43_571 ();
 sg13g2_fill_1 FILLER_43_575 ();
 sg13g2_decap_4 FILLER_43_586 ();
 sg13g2_fill_1 FILLER_43_590 ();
 sg13g2_decap_8 FILLER_43_596 ();
 sg13g2_decap_4 FILLER_43_603 ();
 sg13g2_fill_1 FILLER_43_607 ();
 sg13g2_fill_1 FILLER_43_613 ();
 sg13g2_decap_4 FILLER_43_627 ();
 sg13g2_decap_8 FILLER_43_715 ();
 sg13g2_decap_8 FILLER_43_722 ();
 sg13g2_decap_8 FILLER_43_729 ();
 sg13g2_decap_4 FILLER_43_749 ();
 sg13g2_decap_4 FILLER_43_766 ();
 sg13g2_fill_2 FILLER_43_770 ();
 sg13g2_fill_2 FILLER_43_790 ();
 sg13g2_fill_2 FILLER_43_797 ();
 sg13g2_decap_8 FILLER_43_831 ();
 sg13g2_decap_4 FILLER_43_838 ();
 sg13g2_fill_2 FILLER_43_842 ();
 sg13g2_decap_4 FILLER_43_849 ();
 sg13g2_fill_1 FILLER_43_853 ();
 sg13g2_fill_2 FILLER_43_860 ();
 sg13g2_fill_2 FILLER_43_917 ();
 sg13g2_fill_2 FILLER_43_945 ();
 sg13g2_fill_2 FILLER_43_981 ();
 sg13g2_fill_1 FILLER_43_983 ();
 sg13g2_fill_2 FILLER_43_989 ();
 sg13g2_fill_1 FILLER_43_991 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_fill_2 FILLER_44_56 ();
 sg13g2_fill_2 FILLER_44_71 ();
 sg13g2_decap_8 FILLER_44_83 ();
 sg13g2_decap_4 FILLER_44_94 ();
 sg13g2_decap_4 FILLER_44_107 ();
 sg13g2_decap_4 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_149 ();
 sg13g2_decap_4 FILLER_44_156 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_183 ();
 sg13g2_fill_1 FILLER_44_185 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_237 ();
 sg13g2_fill_1 FILLER_44_255 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_fill_1 FILLER_44_280 ();
 sg13g2_decap_4 FILLER_44_323 ();
 sg13g2_fill_2 FILLER_44_338 ();
 sg13g2_decap_4 FILLER_44_369 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_404 ();
 sg13g2_fill_2 FILLER_44_463 ();
 sg13g2_fill_2 FILLER_44_492 ();
 sg13g2_fill_1 FILLER_44_494 ();
 sg13g2_fill_2 FILLER_44_501 ();
 sg13g2_fill_1 FILLER_44_503 ();
 sg13g2_fill_2 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_562 ();
 sg13g2_decap_8 FILLER_44_569 ();
 sg13g2_fill_2 FILLER_44_589 ();
 sg13g2_decap_4 FILLER_44_618 ();
 sg13g2_fill_2 FILLER_44_622 ();
 sg13g2_fill_1 FILLER_44_645 ();
 sg13g2_fill_2 FILLER_44_673 ();
 sg13g2_fill_1 FILLER_44_675 ();
 sg13g2_fill_2 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_703 ();
 sg13g2_fill_2 FILLER_44_713 ();
 sg13g2_decap_8 FILLER_44_748 ();
 sg13g2_decap_4 FILLER_44_755 ();
 sg13g2_fill_1 FILLER_44_785 ();
 sg13g2_fill_2 FILLER_44_805 ();
 sg13g2_fill_1 FILLER_44_807 ();
 sg13g2_decap_8 FILLER_44_890 ();
 sg13g2_decap_4 FILLER_44_897 ();
 sg13g2_fill_2 FILLER_44_901 ();
 sg13g2_decap_8 FILLER_44_943 ();
 sg13g2_fill_2 FILLER_44_1027 ();
 sg13g2_fill_2 FILLER_45_46 ();
 sg13g2_decap_4 FILLER_45_150 ();
 sg13g2_fill_2 FILLER_45_154 ();
 sg13g2_decap_4 FILLER_45_192 ();
 sg13g2_fill_1 FILLER_45_196 ();
 sg13g2_decap_4 FILLER_45_216 ();
 sg13g2_fill_1 FILLER_45_220 ();
 sg13g2_decap_8 FILLER_45_229 ();
 sg13g2_decap_4 FILLER_45_236 ();
 sg13g2_fill_1 FILLER_45_240 ();
 sg13g2_decap_8 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_271 ();
 sg13g2_decap_8 FILLER_45_278 ();
 sg13g2_decap_4 FILLER_45_285 ();
 sg13g2_fill_2 FILLER_45_289 ();
 sg13g2_fill_2 FILLER_45_313 ();
 sg13g2_fill_1 FILLER_45_315 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_decap_8 FILLER_45_328 ();
 sg13g2_decap_4 FILLER_45_335 ();
 sg13g2_fill_1 FILLER_45_339 ();
 sg13g2_decap_4 FILLER_45_362 ();
 sg13g2_fill_2 FILLER_45_366 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_fill_2 FILLER_45_402 ();
 sg13g2_fill_1 FILLER_45_404 ();
 sg13g2_fill_2 FILLER_45_433 ();
 sg13g2_fill_1 FILLER_45_435 ();
 sg13g2_decap_4 FILLER_45_441 ();
 sg13g2_fill_1 FILLER_45_445 ();
 sg13g2_fill_1 FILLER_45_493 ();
 sg13g2_fill_1 FILLER_45_521 ();
 sg13g2_fill_1 FILLER_45_555 ();
 sg13g2_decap_8 FILLER_45_570 ();
 sg13g2_fill_2 FILLER_45_577 ();
 sg13g2_fill_1 FILLER_45_579 ();
 sg13g2_fill_1 FILLER_45_593 ();
 sg13g2_fill_2 FILLER_45_621 ();
 sg13g2_fill_1 FILLER_45_623 ();
 sg13g2_fill_2 FILLER_45_645 ();
 sg13g2_fill_1 FILLER_45_647 ();
 sg13g2_fill_2 FILLER_45_662 ();
 sg13g2_fill_2 FILLER_45_677 ();
 sg13g2_decap_8 FILLER_45_706 ();
 sg13g2_decap_4 FILLER_45_728 ();
 sg13g2_decap_4 FILLER_45_759 ();
 sg13g2_fill_1 FILLER_45_763 ();
 sg13g2_fill_2 FILLER_45_815 ();
 sg13g2_fill_2 FILLER_45_841 ();
 sg13g2_fill_1 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_849 ();
 sg13g2_fill_1 FILLER_45_862 ();
 sg13g2_fill_2 FILLER_45_880 ();
 sg13g2_fill_1 FILLER_45_882 ();
 sg13g2_fill_2 FILLER_45_902 ();
 sg13g2_fill_1 FILLER_45_904 ();
 sg13g2_fill_1 FILLER_45_938 ();
 sg13g2_decap_4 FILLER_45_966 ();
 sg13g2_fill_1 FILLER_45_970 ();
 sg13g2_decap_8 FILLER_45_988 ();
 sg13g2_decap_8 FILLER_45_1013 ();
 sg13g2_decap_8 FILLER_45_1020 ();
 sg13g2_fill_2 FILLER_45_1027 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_2 FILLER_46_36 ();
 sg13g2_fill_1 FILLER_46_69 ();
 sg13g2_decap_4 FILLER_46_97 ();
 sg13g2_fill_1 FILLER_46_101 ();
 sg13g2_decap_8 FILLER_46_145 ();
 sg13g2_decap_8 FILLER_46_152 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_161 ();
 sg13g2_fill_1 FILLER_46_176 ();
 sg13g2_decap_8 FILLER_46_185 ();
 sg13g2_decap_8 FILLER_46_192 ();
 sg13g2_decap_4 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_208 ();
 sg13g2_fill_2 FILLER_46_215 ();
 sg13g2_fill_2 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_fill_1 FILLER_46_287 ();
 sg13g2_decap_4 FILLER_46_334 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_350 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_1 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_447 ();
 sg13g2_decap_8 FILLER_46_454 ();
 sg13g2_fill_2 FILLER_46_461 ();
 sg13g2_fill_1 FILLER_46_471 ();
 sg13g2_decap_4 FILLER_46_534 ();
 sg13g2_decap_8 FILLER_46_571 ();
 sg13g2_decap_8 FILLER_46_578 ();
 sg13g2_fill_2 FILLER_46_585 ();
 sg13g2_fill_1 FILLER_46_587 ();
 sg13g2_decap_4 FILLER_46_627 ();
 sg13g2_decap_4 FILLER_46_648 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_fill_2 FILLER_46_664 ();
 sg13g2_decap_4 FILLER_46_698 ();
 sg13g2_fill_1 FILLER_46_702 ();
 sg13g2_fill_2 FILLER_46_751 ();
 sg13g2_fill_1 FILLER_46_753 ();
 sg13g2_decap_4 FILLER_46_767 ();
 sg13g2_fill_2 FILLER_46_771 ();
 sg13g2_fill_2 FILLER_46_786 ();
 sg13g2_fill_1 FILLER_46_788 ();
 sg13g2_decap_4 FILLER_46_831 ();
 sg13g2_fill_1 FILLER_46_848 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_4 FILLER_46_938 ();
 sg13g2_fill_2 FILLER_46_942 ();
 sg13g2_decap_4 FILLER_46_957 ();
 sg13g2_fill_2 FILLER_46_961 ();
 sg13g2_fill_2 FILLER_46_972 ();
 sg13g2_decap_8 FILLER_46_1016 ();
 sg13g2_decap_4 FILLER_46_1023 ();
 sg13g2_fill_2 FILLER_46_1027 ();
 sg13g2_decap_4 FILLER_47_4 ();
 sg13g2_fill_1 FILLER_47_8 ();
 sg13g2_fill_1 FILLER_47_28 ();
 sg13g2_fill_1 FILLER_47_41 ();
 sg13g2_fill_1 FILLER_47_93 ();
 sg13g2_fill_2 FILLER_47_127 ();
 sg13g2_decap_8 FILLER_47_152 ();
 sg13g2_decap_8 FILLER_47_159 ();
 sg13g2_fill_2 FILLER_47_166 ();
 sg13g2_fill_1 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_179 ();
 sg13g2_decap_4 FILLER_47_186 ();
 sg13g2_decap_4 FILLER_47_216 ();
 sg13g2_fill_1 FILLER_47_220 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_fill_1 FILLER_47_255 ();
 sg13g2_fill_2 FILLER_47_261 ();
 sg13g2_fill_1 FILLER_47_263 ();
 sg13g2_decap_8 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_decap_8 FILLER_47_304 ();
 sg13g2_fill_2 FILLER_47_332 ();
 sg13g2_fill_2 FILLER_47_357 ();
 sg13g2_fill_1 FILLER_47_359 ();
 sg13g2_fill_1 FILLER_47_366 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_2 FILLER_47_414 ();
 sg13g2_fill_1 FILLER_47_416 ();
 sg13g2_decap_8 FILLER_47_475 ();
 sg13g2_decap_8 FILLER_47_482 ();
 sg13g2_decap_4 FILLER_47_489 ();
 sg13g2_fill_1 FILLER_47_493 ();
 sg13g2_fill_2 FILLER_47_509 ();
 sg13g2_decap_4 FILLER_47_538 ();
 sg13g2_decap_4 FILLER_47_587 ();
 sg13g2_fill_2 FILLER_47_596 ();
 sg13g2_fill_2 FILLER_47_640 ();
 sg13g2_fill_1 FILLER_47_642 ();
 sg13g2_decap_4 FILLER_47_648 ();
 sg13g2_fill_2 FILLER_47_652 ();
 sg13g2_decap_4 FILLER_47_659 ();
 sg13g2_fill_1 FILLER_47_663 ();
 sg13g2_fill_2 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_692 ();
 sg13g2_decap_8 FILLER_47_752 ();
 sg13g2_decap_4 FILLER_47_772 ();
 sg13g2_decap_8 FILLER_47_855 ();
 sg13g2_decap_8 FILLER_47_862 ();
 sg13g2_decap_8 FILLER_47_872 ();
 sg13g2_fill_1 FILLER_47_884 ();
 sg13g2_fill_2 FILLER_47_917 ();
 sg13g2_fill_1 FILLER_47_919 ();
 sg13g2_fill_1 FILLER_47_925 ();
 sg13g2_decap_8 FILLER_47_953 ();
 sg13g2_fill_1 FILLER_47_960 ();
 sg13g2_fill_2 FILLER_47_1000 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_1 FILLER_48_25 ();
 sg13g2_fill_1 FILLER_48_35 ();
 sg13g2_fill_1 FILLER_48_49 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_fill_2 FILLER_48_130 ();
 sg13g2_decap_8 FILLER_48_160 ();
 sg13g2_fill_1 FILLER_48_167 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_decap_4 FILLER_48_232 ();
 sg13g2_fill_1 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_261 ();
 sg13g2_decap_4 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_fill_1 FILLER_48_314 ();
 sg13g2_decap_4 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_373 ();
 sg13g2_fill_2 FILLER_48_387 ();
 sg13g2_decap_8 FILLER_48_398 ();
 sg13g2_decap_8 FILLER_48_405 ();
 sg13g2_decap_8 FILLER_48_412 ();
 sg13g2_decap_8 FILLER_48_419 ();
 sg13g2_fill_2 FILLER_48_426 ();
 sg13g2_fill_1 FILLER_48_428 ();
 sg13g2_fill_2 FILLER_48_443 ();
 sg13g2_fill_1 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_484 ();
 sg13g2_decap_4 FILLER_48_491 ();
 sg13g2_fill_2 FILLER_48_495 ();
 sg13g2_decap_8 FILLER_48_513 ();
 sg13g2_fill_2 FILLER_48_520 ();
 sg13g2_decap_8 FILLER_48_531 ();
 sg13g2_fill_1 FILLER_48_538 ();
 sg13g2_decap_8 FILLER_48_565 ();
 sg13g2_decap_8 FILLER_48_572 ();
 sg13g2_decap_4 FILLER_48_579 ();
 sg13g2_fill_1 FILLER_48_583 ();
 sg13g2_fill_2 FILLER_48_642 ();
 sg13g2_fill_2 FILLER_48_649 ();
 sg13g2_fill_2 FILLER_48_661 ();
 sg13g2_fill_1 FILLER_48_663 ();
 sg13g2_fill_1 FILLER_48_726 ();
 sg13g2_fill_2 FILLER_48_758 ();
 sg13g2_fill_1 FILLER_48_760 ();
 sg13g2_fill_2 FILLER_48_809 ();
 sg13g2_decap_8 FILLER_48_814 ();
 sg13g2_fill_2 FILLER_48_883 ();
 sg13g2_decap_4 FILLER_48_906 ();
 sg13g2_decap_4 FILLER_48_946 ();
 sg13g2_fill_2 FILLER_48_950 ();
 sg13g2_fill_2 FILLER_48_958 ();
 sg13g2_fill_2 FILLER_48_981 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_89 ();
 sg13g2_fill_2 FILLER_49_101 ();
 sg13g2_fill_2 FILLER_49_113 ();
 sg13g2_fill_1 FILLER_49_115 ();
 sg13g2_decap_4 FILLER_49_129 ();
 sg13g2_decap_4 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_fill_1 FILLER_49_224 ();
 sg13g2_decap_4 FILLER_49_255 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_fill_2 FILLER_49_301 ();
 sg13g2_fill_2 FILLER_49_312 ();
 sg13g2_fill_1 FILLER_49_314 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_fill_1 FILLER_49_324 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_fill_1 FILLER_49_350 ();
 sg13g2_fill_1 FILLER_49_355 ();
 sg13g2_fill_2 FILLER_49_390 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_401 ();
 sg13g2_decap_8 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_4 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_426 ();
 sg13g2_decap_4 FILLER_49_431 ();
 sg13g2_fill_2 FILLER_49_435 ();
 sg13g2_decap_8 FILLER_49_468 ();
 sg13g2_decap_8 FILLER_49_475 ();
 sg13g2_fill_2 FILLER_49_482 ();
 sg13g2_fill_2 FILLER_49_497 ();
 sg13g2_fill_1 FILLER_49_505 ();
 sg13g2_fill_2 FILLER_49_515 ();
 sg13g2_fill_2 FILLER_49_535 ();
 sg13g2_fill_1 FILLER_49_537 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_decap_4 FILLER_49_571 ();
 sg13g2_fill_1 FILLER_49_575 ();
 sg13g2_decap_4 FILLER_49_608 ();
 sg13g2_fill_2 FILLER_49_668 ();
 sg13g2_fill_1 FILLER_49_670 ();
 sg13g2_fill_2 FILLER_49_713 ();
 sg13g2_fill_2 FILLER_49_731 ();
 sg13g2_fill_1 FILLER_49_745 ();
 sg13g2_decap_8 FILLER_49_752 ();
 sg13g2_fill_2 FILLER_49_759 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_786 ();
 sg13g2_fill_2 FILLER_49_793 ();
 sg13g2_decap_8 FILLER_49_801 ();
 sg13g2_decap_4 FILLER_49_808 ();
 sg13g2_fill_1 FILLER_49_821 ();
 sg13g2_decap_8 FILLER_49_832 ();
 sg13g2_fill_2 FILLER_49_839 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_4 FILLER_49_863 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_888 ();
 sg13g2_decap_8 FILLER_49_895 ();
 sg13g2_decap_4 FILLER_49_902 ();
 sg13g2_fill_2 FILLER_49_906 ();
 sg13g2_fill_2 FILLER_49_946 ();
 sg13g2_fill_1 FILLER_49_948 ();
 sg13g2_decap_4 FILLER_49_954 ();
 sg13g2_fill_2 FILLER_49_958 ();
 sg13g2_fill_1 FILLER_49_965 ();
 sg13g2_decap_8 FILLER_49_970 ();
 sg13g2_fill_1 FILLER_49_977 ();
 sg13g2_decap_4 FILLER_49_987 ();
 sg13g2_fill_1 FILLER_49_991 ();
 sg13g2_fill_1 FILLER_49_1001 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_fill_1 FILLER_50_76 ();
 sg13g2_fill_1 FILLER_50_86 ();
 sg13g2_fill_2 FILLER_50_142 ();
 sg13g2_fill_2 FILLER_50_153 ();
 sg13g2_fill_1 FILLER_50_155 ();
 sg13g2_decap_8 FILLER_50_247 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_decap_8 FILLER_50_285 ();
 sg13g2_decap_4 FILLER_50_292 ();
 sg13g2_fill_2 FILLER_50_296 ();
 sg13g2_decap_4 FILLER_50_303 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_decap_8 FILLER_50_334 ();
 sg13g2_decap_4 FILLER_50_341 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_2 FILLER_50_378 ();
 sg13g2_fill_1 FILLER_50_380 ();
 sg13g2_fill_2 FILLER_50_410 ();
 sg13g2_fill_1 FILLER_50_422 ();
 sg13g2_fill_1 FILLER_50_439 ();
 sg13g2_decap_4 FILLER_50_451 ();
 sg13g2_decap_8 FILLER_50_464 ();
 sg13g2_decap_8 FILLER_50_471 ();
 sg13g2_decap_8 FILLER_50_478 ();
 sg13g2_decap_4 FILLER_50_512 ();
 sg13g2_fill_1 FILLER_50_516 ();
 sg13g2_decap_8 FILLER_50_558 ();
 sg13g2_fill_2 FILLER_50_602 ();
 sg13g2_fill_1 FILLER_50_604 ();
 sg13g2_decap_8 FILLER_50_631 ();
 sg13g2_fill_2 FILLER_50_638 ();
 sg13g2_decap_8 FILLER_50_697 ();
 sg13g2_decap_4 FILLER_50_704 ();
 sg13g2_fill_1 FILLER_50_708 ();
 sg13g2_fill_2 FILLER_50_727 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_fill_1 FILLER_50_767 ();
 sg13g2_fill_2 FILLER_50_795 ();
 sg13g2_fill_1 FILLER_50_797 ();
 sg13g2_decap_8 FILLER_50_832 ();
 sg13g2_decap_4 FILLER_50_839 ();
 sg13g2_fill_1 FILLER_50_843 ();
 sg13g2_decap_8 FILLER_50_857 ();
 sg13g2_decap_4 FILLER_50_864 ();
 sg13g2_fill_2 FILLER_50_868 ();
 sg13g2_decap_4 FILLER_50_879 ();
 sg13g2_decap_4 FILLER_50_904 ();
 sg13g2_fill_2 FILLER_50_911 ();
 sg13g2_fill_1 FILLER_50_913 ();
 sg13g2_fill_1 FILLER_50_927 ();
 sg13g2_fill_2 FILLER_50_943 ();
 sg13g2_fill_1 FILLER_50_989 ();
 sg13g2_decap_8 FILLER_50_1018 ();
 sg13g2_decap_4 FILLER_50_1025 ();
 sg13g2_fill_2 FILLER_51_77 ();
 sg13g2_fill_1 FILLER_51_79 ();
 sg13g2_fill_2 FILLER_51_104 ();
 sg13g2_fill_1 FILLER_51_106 ();
 sg13g2_fill_2 FILLER_51_116 ();
 sg13g2_fill_1 FILLER_51_118 ();
 sg13g2_decap_8 FILLER_51_128 ();
 sg13g2_decap_4 FILLER_51_135 ();
 sg13g2_fill_2 FILLER_51_139 ();
 sg13g2_fill_2 FILLER_51_168 ();
 sg13g2_fill_1 FILLER_51_170 ();
 sg13g2_fill_2 FILLER_51_200 ();
 sg13g2_fill_2 FILLER_51_212 ();
 sg13g2_fill_2 FILLER_51_233 ();
 sg13g2_decap_8 FILLER_51_248 ();
 sg13g2_decap_4 FILLER_51_255 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_277 ();
 sg13g2_fill_2 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_358 ();
 sg13g2_fill_1 FILLER_51_360 ();
 sg13g2_fill_2 FILLER_51_387 ();
 sg13g2_decap_8 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_410 ();
 sg13g2_fill_2 FILLER_51_448 ();
 sg13g2_fill_1 FILLER_51_450 ();
 sg13g2_fill_2 FILLER_51_469 ();
 sg13g2_decap_4 FILLER_51_487 ();
 sg13g2_decap_4 FILLER_51_501 ();
 sg13g2_fill_1 FILLER_51_505 ();
 sg13g2_fill_1 FILLER_51_519 ();
 sg13g2_decap_4 FILLER_51_526 ();
 sg13g2_decap_4 FILLER_51_563 ();
 sg13g2_fill_2 FILLER_51_567 ();
 sg13g2_fill_1 FILLER_51_584 ();
 sg13g2_fill_1 FILLER_51_603 ();
 sg13g2_fill_1 FILLER_51_610 ();
 sg13g2_fill_2 FILLER_51_651 ();
 sg13g2_fill_1 FILLER_51_653 ();
 sg13g2_decap_8 FILLER_51_658 ();
 sg13g2_decap_4 FILLER_51_665 ();
 sg13g2_fill_2 FILLER_51_711 ();
 sg13g2_fill_1 FILLER_51_713 ();
 sg13g2_decap_8 FILLER_51_737 ();
 sg13g2_decap_8 FILLER_51_744 ();
 sg13g2_fill_1 FILLER_51_751 ();
 sg13g2_fill_1 FILLER_51_792 ();
 sg13g2_fill_2 FILLER_51_825 ();
 sg13g2_fill_2 FILLER_51_889 ();
 sg13g2_fill_2 FILLER_51_923 ();
 sg13g2_fill_1 FILLER_51_925 ();
 sg13g2_decap_8 FILLER_51_967 ();
 sg13g2_fill_1 FILLER_52_51 ();
 sg13g2_decap_4 FILLER_52_133 ();
 sg13g2_decap_4 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_194 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_222 ();
 sg13g2_decap_8 FILLER_52_229 ();
 sg13g2_decap_4 FILLER_52_236 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_decap_8 FILLER_52_247 ();
 sg13g2_decap_8 FILLER_52_254 ();
 sg13g2_decap_4 FILLER_52_261 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_4 FILLER_52_280 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_decap_8 FILLER_52_340 ();
 sg13g2_fill_1 FILLER_52_347 ();
 sg13g2_decap_4 FILLER_52_375 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_4 FILLER_52_392 ();
 sg13g2_fill_1 FILLER_52_396 ();
 sg13g2_fill_1 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_decap_8 FILLER_52_415 ();
 sg13g2_decap_4 FILLER_52_422 ();
 sg13g2_fill_2 FILLER_52_426 ();
 sg13g2_fill_2 FILLER_52_437 ();
 sg13g2_fill_1 FILLER_52_444 ();
 sg13g2_fill_1 FILLER_52_450 ();
 sg13g2_decap_8 FILLER_52_500 ();
 sg13g2_fill_1 FILLER_52_507 ();
 sg13g2_fill_2 FILLER_52_540 ();
 sg13g2_fill_1 FILLER_52_542 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_decap_8 FILLER_52_562 ();
 sg13g2_fill_2 FILLER_52_569 ();
 sg13g2_fill_1 FILLER_52_571 ();
 sg13g2_fill_1 FILLER_52_606 ();
 sg13g2_decap_8 FILLER_52_612 ();
 sg13g2_decap_4 FILLER_52_619 ();
 sg13g2_decap_8 FILLER_52_632 ();
 sg13g2_decap_8 FILLER_52_639 ();
 sg13g2_decap_8 FILLER_52_646 ();
 sg13g2_decap_4 FILLER_52_653 ();
 sg13g2_fill_2 FILLER_52_657 ();
 sg13g2_decap_4 FILLER_52_665 ();
 sg13g2_decap_4 FILLER_52_678 ();
 sg13g2_fill_1 FILLER_52_682 ();
 sg13g2_fill_1 FILLER_52_748 ();
 sg13g2_fill_2 FILLER_52_762 ();
 sg13g2_decap_4 FILLER_52_791 ();
 sg13g2_fill_1 FILLER_52_795 ();
 sg13g2_decap_8 FILLER_52_829 ();
 sg13g2_fill_2 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_838 ();
 sg13g2_fill_1 FILLER_52_848 ();
 sg13g2_fill_2 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_862 ();
 sg13g2_fill_2 FILLER_52_869 ();
 sg13g2_decap_4 FILLER_52_897 ();
 sg13g2_decap_4 FILLER_52_906 ();
 sg13g2_fill_2 FILLER_52_910 ();
 sg13g2_decap_8 FILLER_52_935 ();
 sg13g2_decap_8 FILLER_52_942 ();
 sg13g2_fill_2 FILLER_52_949 ();
 sg13g2_decap_4 FILLER_52_968 ();
 sg13g2_fill_2 FILLER_52_972 ();
 sg13g2_fill_2 FILLER_52_1026 ();
 sg13g2_fill_1 FILLER_52_1028 ();
 sg13g2_decap_4 FILLER_53_4 ();
 sg13g2_fill_2 FILLER_53_8 ();
 sg13g2_decap_8 FILLER_53_38 ();
 sg13g2_decap_4 FILLER_53_45 ();
 sg13g2_fill_2 FILLER_53_49 ();
 sg13g2_decap_4 FILLER_53_55 ();
 sg13g2_fill_2 FILLER_53_94 ();
 sg13g2_fill_1 FILLER_53_96 ();
 sg13g2_decap_8 FILLER_53_114 ();
 sg13g2_decap_4 FILLER_53_121 ();
 sg13g2_fill_2 FILLER_53_125 ();
 sg13g2_fill_2 FILLER_53_146 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_decap_8 FILLER_53_159 ();
 sg13g2_fill_2 FILLER_53_226 ();
 sg13g2_fill_2 FILLER_53_254 ();
 sg13g2_fill_2 FILLER_53_263 ();
 sg13g2_decap_4 FILLER_53_273 ();
 sg13g2_decap_4 FILLER_53_308 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_decap_8 FILLER_53_358 ();
 sg13g2_decap_8 FILLER_53_365 ();
 sg13g2_fill_2 FILLER_53_372 ();
 sg13g2_fill_1 FILLER_53_374 ();
 sg13g2_decap_4 FILLER_53_401 ();
 sg13g2_fill_2 FILLER_53_405 ();
 sg13g2_fill_2 FILLER_53_434 ();
 sg13g2_fill_1 FILLER_53_436 ();
 sg13g2_fill_2 FILLER_53_449 ();
 sg13g2_decap_4 FILLER_53_469 ();
 sg13g2_decap_8 FILLER_53_505 ();
 sg13g2_fill_1 FILLER_53_512 ();
 sg13g2_fill_1 FILLER_53_526 ();
 sg13g2_fill_1 FILLER_53_547 ();
 sg13g2_fill_2 FILLER_53_561 ();
 sg13g2_fill_1 FILLER_53_563 ();
 sg13g2_fill_2 FILLER_53_577 ();
 sg13g2_fill_1 FILLER_53_579 ();
 sg13g2_fill_1 FILLER_53_585 ();
 sg13g2_decap_8 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_614 ();
 sg13g2_fill_2 FILLER_53_621 ();
 sg13g2_fill_1 FILLER_53_623 ();
 sg13g2_fill_1 FILLER_53_645 ();
 sg13g2_decap_8 FILLER_53_678 ();
 sg13g2_fill_1 FILLER_53_685 ();
 sg13g2_fill_1 FILLER_53_712 ();
 sg13g2_fill_1 FILLER_53_750 ();
 sg13g2_decap_8 FILLER_53_764 ();
 sg13g2_fill_2 FILLER_53_771 ();
 sg13g2_fill_1 FILLER_53_773 ();
 sg13g2_fill_2 FILLER_53_795 ();
 sg13g2_fill_1 FILLER_53_797 ();
 sg13g2_fill_1 FILLER_53_803 ();
 sg13g2_fill_2 FILLER_53_829 ();
 sg13g2_decap_8 FILLER_53_842 ();
 sg13g2_fill_1 FILLER_53_864 ();
 sg13g2_decap_4 FILLER_53_889 ();
 sg13g2_decap_4 FILLER_53_901 ();
 sg13g2_fill_2 FILLER_53_905 ();
 sg13g2_fill_2 FILLER_53_920 ();
 sg13g2_fill_1 FILLER_53_922 ();
 sg13g2_decap_8 FILLER_53_936 ();
 sg13g2_decap_4 FILLER_53_943 ();
 sg13g2_decap_4 FILLER_53_975 ();
 sg13g2_fill_1 FILLER_53_979 ();
 sg13g2_fill_2 FILLER_53_985 ();
 sg13g2_fill_1 FILLER_53_987 ();
 sg13g2_decap_4 FILLER_53_1024 ();
 sg13g2_fill_1 FILLER_53_1028 ();
 sg13g2_decap_4 FILLER_54_37 ();
 sg13g2_decap_4 FILLER_54_54 ();
 sg13g2_fill_1 FILLER_54_58 ();
 sg13g2_fill_1 FILLER_54_117 ();
 sg13g2_fill_2 FILLER_54_213 ();
 sg13g2_decap_4 FILLER_54_219 ();
 sg13g2_fill_2 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_4 FILLER_54_258 ();
 sg13g2_fill_1 FILLER_54_267 ();
 sg13g2_decap_8 FILLER_54_274 ();
 sg13g2_decap_8 FILLER_54_281 ();
 sg13g2_decap_8 FILLER_54_288 ();
 sg13g2_decap_8 FILLER_54_295 ();
 sg13g2_decap_4 FILLER_54_340 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_2 FILLER_54_441 ();
 sg13g2_fill_2 FILLER_54_447 ();
 sg13g2_fill_1 FILLER_54_463 ();
 sg13g2_decap_4 FILLER_54_520 ();
 sg13g2_fill_2 FILLER_54_524 ();
 sg13g2_fill_2 FILLER_54_562 ();
 sg13g2_decap_4 FILLER_54_599 ();
 sg13g2_decap_4 FILLER_54_651 ();
 sg13g2_fill_1 FILLER_54_688 ();
 sg13g2_fill_2 FILLER_54_729 ();
 sg13g2_fill_2 FILLER_54_759 ();
 sg13g2_fill_1 FILLER_54_788 ();
 sg13g2_decap_4 FILLER_54_827 ();
 sg13g2_fill_1 FILLER_54_831 ();
 sg13g2_fill_1 FILLER_54_870 ();
 sg13g2_decap_4 FILLER_54_919 ();
 sg13g2_fill_1 FILLER_54_923 ();
 sg13g2_fill_2 FILLER_54_964 ();
 sg13g2_fill_1 FILLER_54_966 ();
 sg13g2_fill_2 FILLER_54_992 ();
 sg13g2_decap_8 FILLER_54_1021 ();
 sg13g2_fill_1 FILLER_54_1028 ();
 sg13g2_decap_8 FILLER_55_4 ();
 sg13g2_decap_4 FILLER_55_11 ();
 sg13g2_fill_2 FILLER_55_15 ();
 sg13g2_fill_2 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_206 ();
 sg13g2_decap_8 FILLER_55_213 ();
 sg13g2_decap_4 FILLER_55_220 ();
 sg13g2_decap_4 FILLER_55_238 ();
 sg13g2_decap_4 FILLER_55_258 ();
 sg13g2_fill_2 FILLER_55_270 ();
 sg13g2_decap_8 FILLER_55_312 ();
 sg13g2_decap_4 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_332 ();
 sg13g2_decap_4 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_342 ();
 sg13g2_decap_4 FILLER_55_351 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_374 ();
 sg13g2_fill_1 FILLER_55_376 ();
 sg13g2_decap_4 FILLER_55_404 ();
 sg13g2_fill_2 FILLER_55_417 ();
 sg13g2_fill_1 FILLER_55_419 ();
 sg13g2_decap_8 FILLER_55_446 ();
 sg13g2_decap_8 FILLER_55_453 ();
 sg13g2_decap_8 FILLER_55_464 ();
 sg13g2_decap_8 FILLER_55_471 ();
 sg13g2_decap_4 FILLER_55_478 ();
 sg13g2_fill_1 FILLER_55_482 ();
 sg13g2_decap_4 FILLER_55_488 ();
 sg13g2_fill_1 FILLER_55_492 ();
 sg13g2_fill_2 FILLER_55_504 ();
 sg13g2_fill_1 FILLER_55_506 ();
 sg13g2_fill_2 FILLER_55_544 ();
 sg13g2_decap_4 FILLER_55_569 ();
 sg13g2_fill_1 FILLER_55_573 ();
 sg13g2_decap_4 FILLER_55_583 ();
 sg13g2_fill_1 FILLER_55_587 ();
 sg13g2_decap_8 FILLER_55_596 ();
 sg13g2_decap_8 FILLER_55_603 ();
 sg13g2_decap_8 FILLER_55_610 ();
 sg13g2_fill_2 FILLER_55_654 ();
 sg13g2_fill_2 FILLER_55_661 ();
 sg13g2_fill_1 FILLER_55_676 ();
 sg13g2_decap_8 FILLER_55_692 ();
 sg13g2_decap_4 FILLER_55_699 ();
 sg13g2_fill_2 FILLER_55_729 ();
 sg13g2_fill_1 FILLER_55_731 ();
 sg13g2_fill_2 FILLER_55_741 ();
 sg13g2_decap_4 FILLER_55_765 ();
 sg13g2_fill_2 FILLER_55_789 ();
 sg13g2_fill_1 FILLER_55_791 ();
 sg13g2_fill_1 FILLER_55_797 ();
 sg13g2_fill_1 FILLER_55_815 ();
 sg13g2_decap_4 FILLER_55_822 ();
 sg13g2_fill_2 FILLER_55_858 ();
 sg13g2_fill_1 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_55_883 ();
 sg13g2_decap_8 FILLER_55_940 ();
 sg13g2_decap_8 FILLER_55_947 ();
 sg13g2_decap_8 FILLER_55_988 ();
 sg13g2_decap_8 FILLER_55_1013 ();
 sg13g2_decap_8 FILLER_55_1020 ();
 sg13g2_fill_2 FILLER_55_1027 ();
 sg13g2_fill_2 FILLER_56_40 ();
 sg13g2_fill_1 FILLER_56_42 ();
 sg13g2_decap_4 FILLER_56_75 ();
 sg13g2_decap_4 FILLER_56_111 ();
 sg13g2_fill_2 FILLER_56_146 ();
 sg13g2_decap_4 FILLER_56_157 ();
 sg13g2_fill_1 FILLER_56_161 ();
 sg13g2_fill_2 FILLER_56_208 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_2 FILLER_56_230 ();
 sg13g2_fill_1 FILLER_56_232 ();
 sg13g2_fill_2 FILLER_56_251 ();
 sg13g2_fill_2 FILLER_56_261 ();
 sg13g2_fill_1 FILLER_56_263 ();
 sg13g2_decap_4 FILLER_56_269 ();
 sg13g2_decap_4 FILLER_56_286 ();
 sg13g2_fill_2 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_322 ();
 sg13g2_decap_4 FILLER_56_418 ();
 sg13g2_fill_2 FILLER_56_422 ();
 sg13g2_decap_4 FILLER_56_437 ();
 sg13g2_decap_4 FILLER_56_454 ();
 sg13g2_decap_8 FILLER_56_509 ();
 sg13g2_fill_2 FILLER_56_516 ();
 sg13g2_fill_1 FILLER_56_518 ();
 sg13g2_decap_4 FILLER_56_525 ();
 sg13g2_fill_2 FILLER_56_529 ();
 sg13g2_fill_2 FILLER_56_559 ();
 sg13g2_fill_1 FILLER_56_561 ();
 sg13g2_fill_1 FILLER_56_567 ();
 sg13g2_fill_2 FILLER_56_574 ();
 sg13g2_fill_1 FILLER_56_576 ();
 sg13g2_decap_4 FILLER_56_592 ();
 sg13g2_fill_2 FILLER_56_596 ();
 sg13g2_decap_8 FILLER_56_646 ();
 sg13g2_decap_8 FILLER_56_653 ();
 sg13g2_decap_4 FILLER_56_660 ();
 sg13g2_fill_2 FILLER_56_664 ();
 sg13g2_fill_2 FILLER_56_702 ();
 sg13g2_decap_8 FILLER_56_740 ();
 sg13g2_decap_8 FILLER_56_747 ();
 sg13g2_decap_4 FILLER_56_754 ();
 sg13g2_decap_4 FILLER_56_785 ();
 sg13g2_fill_2 FILLER_56_789 ();
 sg13g2_fill_1 FILLER_56_796 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_4 FILLER_56_845 ();
 sg13g2_decap_4 FILLER_56_858 ();
 sg13g2_fill_2 FILLER_56_862 ();
 sg13g2_fill_1 FILLER_56_883 ();
 sg13g2_decap_4 FILLER_56_949 ();
 sg13g2_fill_2 FILLER_56_953 ();
 sg13g2_fill_2 FILLER_56_960 ();
 sg13g2_decap_4 FILLER_56_983 ();
 sg13g2_fill_1 FILLER_56_990 ();
 sg13g2_decap_8 FILLER_56_1018 ();
 sg13g2_decap_4 FILLER_56_1025 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_4 FILLER_57_7 ();
 sg13g2_fill_2 FILLER_57_20 ();
 sg13g2_fill_2 FILLER_57_35 ();
 sg13g2_decap_4 FILLER_57_45 ();
 sg13g2_fill_1 FILLER_57_58 ();
 sg13g2_fill_2 FILLER_57_73 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_4 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_decap_8 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_171 ();
 sg13g2_fill_1 FILLER_57_190 ();
 sg13g2_decap_8 FILLER_57_204 ();
 sg13g2_decap_8 FILLER_57_221 ();
 sg13g2_decap_8 FILLER_57_228 ();
 sg13g2_fill_1 FILLER_57_235 ();
 sg13g2_decap_8 FILLER_57_256 ();
 sg13g2_decap_8 FILLER_57_263 ();
 sg13g2_decap_8 FILLER_57_270 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_decap_8 FILLER_57_282 ();
 sg13g2_decap_8 FILLER_57_289 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_fill_1 FILLER_57_420 ();
 sg13g2_fill_2 FILLER_57_432 ();
 sg13g2_fill_1 FILLER_57_434 ();
 sg13g2_fill_2 FILLER_57_454 ();
 sg13g2_fill_2 FILLER_57_483 ();
 sg13g2_decap_4 FILLER_57_519 ();
 sg13g2_decap_8 FILLER_57_552 ();
 sg13g2_decap_4 FILLER_57_600 ();
 sg13g2_fill_1 FILLER_57_604 ();
 sg13g2_decap_4 FILLER_57_632 ();
 sg13g2_fill_2 FILLER_57_675 ();
 sg13g2_fill_1 FILLER_57_693 ();
 sg13g2_fill_2 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_731 ();
 sg13g2_fill_1 FILLER_57_738 ();
 sg13g2_fill_2 FILLER_57_766 ();
 sg13g2_fill_2 FILLER_57_777 ();
 sg13g2_fill_1 FILLER_57_779 ();
 sg13g2_fill_1 FILLER_57_795 ();
 sg13g2_fill_2 FILLER_57_823 ();
 sg13g2_fill_1 FILLER_57_825 ();
 sg13g2_fill_2 FILLER_57_869 ();
 sg13g2_decap_8 FILLER_57_878 ();
 sg13g2_decap_8 FILLER_57_885 ();
 sg13g2_fill_1 FILLER_57_892 ();
 sg13g2_decap_4 FILLER_57_896 ();
 sg13g2_fill_2 FILLER_57_900 ();
 sg13g2_fill_1 FILLER_57_915 ();
 sg13g2_fill_2 FILLER_57_943 ();
 sg13g2_decap_4 FILLER_57_958 ();
 sg13g2_fill_1 FILLER_57_962 ();
 sg13g2_fill_1 FILLER_57_980 ();
 sg13g2_decap_8 FILLER_57_1017 ();
 sg13g2_decap_4 FILLER_57_1024 ();
 sg13g2_fill_1 FILLER_57_1028 ();
 sg13g2_decap_8 FILLER_58_4 ();
 sg13g2_decap_8 FILLER_58_11 ();
 sg13g2_fill_2 FILLER_58_18 ();
 sg13g2_fill_1 FILLER_58_20 ();
 sg13g2_fill_2 FILLER_58_85 ();
 sg13g2_fill_1 FILLER_58_87 ();
 sg13g2_fill_1 FILLER_58_99 ();
 sg13g2_decap_8 FILLER_58_166 ();
 sg13g2_decap_8 FILLER_58_173 ();
 sg13g2_decap_4 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_200 ();
 sg13g2_decap_4 FILLER_58_206 ();
 sg13g2_decap_8 FILLER_58_214 ();
 sg13g2_decap_8 FILLER_58_253 ();
 sg13g2_decap_8 FILLER_58_260 ();
 sg13g2_decap_4 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_decap_4 FILLER_58_300 ();
 sg13g2_fill_2 FILLER_58_304 ();
 sg13g2_decap_8 FILLER_58_319 ();
 sg13g2_fill_1 FILLER_58_339 ();
 sg13g2_fill_2 FILLER_58_362 ();
 sg13g2_fill_1 FILLER_58_406 ();
 sg13g2_decap_4 FILLER_58_463 ();
 sg13g2_fill_1 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_481 ();
 sg13g2_decap_4 FILLER_58_506 ();
 sg13g2_decap_8 FILLER_58_554 ();
 sg13g2_decap_8 FILLER_58_561 ();
 sg13g2_decap_4 FILLER_58_568 ();
 sg13g2_fill_1 FILLER_58_572 ();
 sg13g2_decap_4 FILLER_58_603 ();
 sg13g2_fill_1 FILLER_58_607 ();
 sg13g2_decap_8 FILLER_58_621 ();
 sg13g2_decap_8 FILLER_58_647 ();
 sg13g2_decap_4 FILLER_58_667 ();
 sg13g2_fill_1 FILLER_58_671 ();
 sg13g2_fill_1 FILLER_58_712 ();
 sg13g2_decap_8 FILLER_58_734 ();
 sg13g2_decap_8 FILLER_58_741 ();
 sg13g2_fill_2 FILLER_58_748 ();
 sg13g2_decap_8 FILLER_58_788 ();
 sg13g2_decap_4 FILLER_58_795 ();
 sg13g2_fill_2 FILLER_58_799 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_4 FILLER_58_828 ();
 sg13g2_fill_1 FILLER_58_832 ();
 sg13g2_decap_4 FILLER_58_860 ();
 sg13g2_decap_8 FILLER_58_871 ();
 sg13g2_decap_4 FILLER_58_878 ();
 sg13g2_fill_2 FILLER_58_882 ();
 sg13g2_fill_1 FILLER_58_889 ();
 sg13g2_decap_4 FILLER_58_899 ();
 sg13g2_fill_2 FILLER_58_916 ();
 sg13g2_decap_4 FILLER_58_940 ();
 sg13g2_fill_1 FILLER_58_944 ();
 sg13g2_decap_8 FILLER_58_958 ();
 sg13g2_decap_8 FILLER_58_965 ();
 sg13g2_fill_1 FILLER_58_972 ();
 sg13g2_fill_2 FILLER_59_27 ();
 sg13g2_fill_1 FILLER_59_56 ();
 sg13g2_decap_4 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_fill_1 FILLER_59_140 ();
 sg13g2_fill_2 FILLER_59_178 ();
 sg13g2_fill_1 FILLER_59_180 ();
 sg13g2_decap_4 FILLER_59_229 ();
 sg13g2_fill_2 FILLER_59_233 ();
 sg13g2_decap_8 FILLER_59_244 ();
 sg13g2_decap_4 FILLER_59_268 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_fill_2 FILLER_59_301 ();
 sg13g2_fill_1 FILLER_59_303 ();
 sg13g2_decap_4 FILLER_59_309 ();
 sg13g2_fill_2 FILLER_59_313 ();
 sg13g2_decap_8 FILLER_59_356 ();
 sg13g2_decap_4 FILLER_59_363 ();
 sg13g2_fill_1 FILLER_59_367 ();
 sg13g2_fill_2 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_decap_8 FILLER_59_418 ();
 sg13g2_fill_1 FILLER_59_425 ();
 sg13g2_decap_4 FILLER_59_456 ();
 sg13g2_fill_1 FILLER_59_500 ();
 sg13g2_decap_8 FILLER_59_510 ();
 sg13g2_decap_8 FILLER_59_517 ();
 sg13g2_fill_2 FILLER_59_524 ();
 sg13g2_fill_1 FILLER_59_526 ();
 sg13g2_fill_1 FILLER_59_533 ();
 sg13g2_decap_8 FILLER_59_543 ();
 sg13g2_decap_4 FILLER_59_550 ();
 sg13g2_fill_2 FILLER_59_554 ();
 sg13g2_fill_2 FILLER_59_561 ();
 sg13g2_decap_8 FILLER_59_569 ();
 sg13g2_decap_8 FILLER_59_576 ();
 sg13g2_decap_8 FILLER_59_583 ();
 sg13g2_fill_2 FILLER_59_590 ();
 sg13g2_fill_1 FILLER_59_592 ();
 sg13g2_fill_2 FILLER_59_609 ();
 sg13g2_fill_2 FILLER_59_624 ();
 sg13g2_fill_1 FILLER_59_626 ();
 sg13g2_fill_2 FILLER_59_645 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_decap_8 FILLER_59_689 ();
 sg13g2_decap_8 FILLER_59_696 ();
 sg13g2_fill_1 FILLER_59_713 ();
 sg13g2_fill_1 FILLER_59_723 ();
 sg13g2_fill_2 FILLER_59_730 ();
 sg13g2_fill_1 FILLER_59_732 ();
 sg13g2_fill_2 FILLER_59_742 ();
 sg13g2_fill_1 FILLER_59_744 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_fill_2 FILLER_59_803 ();
 sg13g2_fill_1 FILLER_59_805 ();
 sg13g2_decap_4 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_839 ();
 sg13g2_fill_1 FILLER_59_846 ();
 sg13g2_fill_1 FILLER_59_856 ();
 sg13g2_fill_1 FILLER_59_879 ();
 sg13g2_decap_8 FILLER_59_909 ();
 sg13g2_decap_8 FILLER_59_943 ();
 sg13g2_fill_1 FILLER_59_980 ();
 sg13g2_fill_2 FILLER_59_999 ();
 sg13g2_fill_1 FILLER_59_1001 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_fill_1 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_27 ();
 sg13g2_decap_4 FILLER_60_50 ();
 sg13g2_fill_2 FILLER_60_54 ();
 sg13g2_fill_1 FILLER_60_69 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_fill_1 FILLER_60_136 ();
 sg13g2_fill_2 FILLER_60_159 ();
 sg13g2_decap_8 FILLER_60_170 ();
 sg13g2_decap_8 FILLER_60_177 ();
 sg13g2_decap_4 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_222 ();
 sg13g2_decap_4 FILLER_60_250 ();
 sg13g2_fill_1 FILLER_60_254 ();
 sg13g2_decap_4 FILLER_60_261 ();
 sg13g2_fill_2 FILLER_60_265 ();
 sg13g2_decap_4 FILLER_60_289 ();
 sg13g2_fill_2 FILLER_60_320 ();
 sg13g2_decap_8 FILLER_60_339 ();
 sg13g2_fill_1 FILLER_60_346 ();
 sg13g2_fill_2 FILLER_60_375 ();
 sg13g2_fill_2 FILLER_60_400 ();
 sg13g2_decap_8 FILLER_60_415 ();
 sg13g2_decap_4 FILLER_60_422 ();
 sg13g2_fill_1 FILLER_60_453 ();
 sg13g2_decap_8 FILLER_60_475 ();
 sg13g2_fill_2 FILLER_60_482 ();
 sg13g2_fill_1 FILLER_60_484 ();
 sg13g2_fill_2 FILLER_60_498 ();
 sg13g2_fill_1 FILLER_60_505 ();
 sg13g2_fill_1 FILLER_60_517 ();
 sg13g2_fill_2 FILLER_60_524 ();
 sg13g2_decap_8 FILLER_60_535 ();
 sg13g2_fill_1 FILLER_60_542 ();
 sg13g2_fill_2 FILLER_60_547 ();
 sg13g2_fill_1 FILLER_60_593 ();
 sg13g2_fill_2 FILLER_60_600 ();
 sg13g2_decap_4 FILLER_60_629 ();
 sg13g2_fill_1 FILLER_60_633 ();
 sg13g2_decap_8 FILLER_60_688 ();
 sg13g2_fill_2 FILLER_60_695 ();
 sg13g2_fill_1 FILLER_60_697 ();
 sg13g2_fill_2 FILLER_60_712 ();
 sg13g2_fill_2 FILLER_60_741 ();
 sg13g2_fill_1 FILLER_60_791 ();
 sg13g2_fill_2 FILLER_60_799 ();
 sg13g2_fill_1 FILLER_60_861 ();
 sg13g2_decap_8 FILLER_60_878 ();
 sg13g2_fill_2 FILLER_60_885 ();
 sg13g2_fill_1 FILLER_60_887 ();
 sg13g2_decap_4 FILLER_60_905 ();
 sg13g2_decap_8 FILLER_60_929 ();
 sg13g2_decap_8 FILLER_60_936 ();
 sg13g2_decap_4 FILLER_60_943 ();
 sg13g2_fill_2 FILLER_60_947 ();
 sg13g2_fill_1 FILLER_60_973 ();
 sg13g2_decap_8 FILLER_60_1014 ();
 sg13g2_decap_8 FILLER_60_1021 ();
 sg13g2_fill_1 FILLER_60_1028 ();
 sg13g2_fill_1 FILLER_61_5 ();
 sg13g2_decap_4 FILLER_61_46 ();
 sg13g2_fill_1 FILLER_61_50 ();
 sg13g2_fill_1 FILLER_61_79 ();
 sg13g2_fill_2 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_138 ();
 sg13g2_fill_1 FILLER_61_145 ();
 sg13g2_decap_4 FILLER_61_168 ();
 sg13g2_decap_4 FILLER_61_249 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_fill_1 FILLER_61_298 ();
 sg13g2_decap_8 FILLER_61_387 ();
 sg13g2_decap_4 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_405 ();
 sg13g2_fill_1 FILLER_61_433 ();
 sg13g2_decap_8 FILLER_61_475 ();
 sg13g2_decap_8 FILLER_61_482 ();
 sg13g2_fill_1 FILLER_61_489 ();
 sg13g2_fill_1 FILLER_61_503 ();
 sg13g2_fill_2 FILLER_61_552 ();
 sg13g2_fill_1 FILLER_61_554 ();
 sg13g2_decap_4 FILLER_61_568 ();
 sg13g2_decap_4 FILLER_61_598 ();
 sg13g2_fill_1 FILLER_61_629 ();
 sg13g2_decap_4 FILLER_61_648 ();
 sg13g2_decap_8 FILLER_61_674 ();
 sg13g2_decap_8 FILLER_61_681 ();
 sg13g2_decap_4 FILLER_61_688 ();
 sg13g2_fill_2 FILLER_61_692 ();
 sg13g2_fill_1 FILLER_61_723 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_decap_8 FILLER_61_742 ();
 sg13g2_decap_4 FILLER_61_749 ();
 sg13g2_fill_2 FILLER_61_753 ();
 sg13g2_decap_8 FILLER_61_760 ();
 sg13g2_fill_2 FILLER_61_767 ();
 sg13g2_fill_1 FILLER_61_769 ();
 sg13g2_fill_1 FILLER_61_776 ();
 sg13g2_fill_2 FILLER_61_782 ();
 sg13g2_fill_1 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_fill_1 FILLER_61_802 ();
 sg13g2_fill_1 FILLER_61_813 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_4 FILLER_61_844 ();
 sg13g2_fill_1 FILLER_61_848 ();
 sg13g2_decap_8 FILLER_61_880 ();
 sg13g2_decap_8 FILLER_61_887 ();
 sg13g2_decap_4 FILLER_61_894 ();
 sg13g2_fill_2 FILLER_61_898 ();
 sg13g2_decap_8 FILLER_61_942 ();
 sg13g2_fill_2 FILLER_61_968 ();
 sg13g2_decap_4 FILLER_61_982 ();
 sg13g2_decap_8 FILLER_61_1013 ();
 sg13g2_decap_8 FILLER_61_1020 ();
 sg13g2_fill_2 FILLER_61_1027 ();
 sg13g2_fill_2 FILLER_62_27 ();
 sg13g2_fill_1 FILLER_62_29 ();
 sg13g2_decap_8 FILLER_62_106 ();
 sg13g2_fill_2 FILLER_62_113 ();
 sg13g2_decap_4 FILLER_62_174 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_decap_4 FILLER_62_212 ();
 sg13g2_decap_8 FILLER_62_226 ();
 sg13g2_decap_8 FILLER_62_261 ();
 sg13g2_decap_8 FILLER_62_268 ();
 sg13g2_decap_4 FILLER_62_306 ();
 sg13g2_fill_2 FILLER_62_310 ();
 sg13g2_decap_4 FILLER_62_321 ();
 sg13g2_fill_1 FILLER_62_325 ();
 sg13g2_fill_2 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_341 ();
 sg13g2_fill_1 FILLER_62_393 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_fill_2 FILLER_62_441 ();
 sg13g2_fill_2 FILLER_62_448 ();
 sg13g2_fill_1 FILLER_62_450 ();
 sg13g2_decap_8 FILLER_62_478 ();
 sg13g2_decap_8 FILLER_62_485 ();
 sg13g2_fill_1 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_529 ();
 sg13g2_decap_8 FILLER_62_552 ();
 sg13g2_fill_1 FILLER_62_559 ();
 sg13g2_fill_2 FILLER_62_572 ();
 sg13g2_fill_1 FILLER_62_574 ();
 sg13g2_decap_8 FILLER_62_596 ();
 sg13g2_fill_1 FILLER_62_603 ();
 sg13g2_decap_4 FILLER_62_622 ();
 sg13g2_fill_1 FILLER_62_632 ();
 sg13g2_fill_2 FILLER_62_646 ();
 sg13g2_fill_1 FILLER_62_648 ();
 sg13g2_decap_4 FILLER_62_698 ();
 sg13g2_fill_1 FILLER_62_733 ();
 sg13g2_decap_4 FILLER_62_740 ();
 sg13g2_fill_2 FILLER_62_744 ();
 sg13g2_fill_2 FILLER_62_755 ();
 sg13g2_fill_1 FILLER_62_757 ();
 sg13g2_fill_2 FILLER_62_763 ();
 sg13g2_fill_1 FILLER_62_765 ();
 sg13g2_decap_4 FILLER_62_772 ();
 sg13g2_fill_1 FILLER_62_785 ();
 sg13g2_fill_1 FILLER_62_794 ();
 sg13g2_decap_8 FILLER_62_803 ();
 sg13g2_fill_2 FILLER_62_810 ();
 sg13g2_decap_8 FILLER_62_839 ();
 sg13g2_fill_2 FILLER_62_846 ();
 sg13g2_fill_1 FILLER_62_848 ();
 sg13g2_fill_1 FILLER_62_862 ();
 sg13g2_fill_2 FILLER_62_889 ();
 sg13g2_fill_1 FILLER_62_891 ();
 sg13g2_fill_2 FILLER_62_962 ();
 sg13g2_fill_2 FILLER_62_968 ();
 sg13g2_decap_4 FILLER_62_976 ();
 sg13g2_decap_8 FILLER_62_1021 ();
 sg13g2_fill_1 FILLER_62_1028 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_decap_4 FILLER_63_46 ();
 sg13g2_fill_2 FILLER_63_68 ();
 sg13g2_fill_2 FILLER_63_107 ();
 sg13g2_fill_2 FILLER_63_145 ();
 sg13g2_fill_1 FILLER_63_147 ();
 sg13g2_decap_4 FILLER_63_180 ();
 sg13g2_decap_8 FILLER_63_215 ();
 sg13g2_decap_4 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_271 ();
 sg13g2_fill_2 FILLER_63_286 ();
 sg13g2_decap_4 FILLER_63_298 ();
 sg13g2_fill_2 FILLER_63_302 ();
 sg13g2_fill_1 FILLER_63_332 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_decap_4 FILLER_63_390 ();
 sg13g2_fill_1 FILLER_63_394 ();
 sg13g2_decap_8 FILLER_63_404 ();
 sg13g2_decap_8 FILLER_63_419 ();
 sg13g2_fill_2 FILLER_63_426 ();
 sg13g2_fill_1 FILLER_63_428 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_fill_2 FILLER_63_455 ();
 sg13g2_fill_2 FILLER_63_479 ();
 sg13g2_fill_1 FILLER_63_481 ();
 sg13g2_fill_2 FILLER_63_501 ();
 sg13g2_fill_1 FILLER_63_503 ();
 sg13g2_fill_2 FILLER_63_559 ();
 sg13g2_fill_1 FILLER_63_561 ();
 sg13g2_decap_4 FILLER_63_598 ();
 sg13g2_fill_1 FILLER_63_602 ();
 sg13g2_fill_2 FILLER_63_621 ();
 sg13g2_fill_1 FILLER_63_645 ();
 sg13g2_decap_4 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_682 ();
 sg13g2_fill_1 FILLER_63_689 ();
 sg13g2_fill_2 FILLER_63_716 ();
 sg13g2_fill_2 FILLER_63_725 ();
 sg13g2_fill_1 FILLER_63_727 ();
 sg13g2_decap_8 FILLER_63_813 ();
 sg13g2_decap_8 FILLER_63_820 ();
 sg13g2_decap_8 FILLER_63_827 ();
 sg13g2_decap_4 FILLER_63_834 ();
 sg13g2_decap_8 FILLER_63_843 ();
 sg13g2_fill_2 FILLER_63_850 ();
 sg13g2_fill_1 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_2 FILLER_63_884 ();
 sg13g2_decap_8 FILLER_63_895 ();
 sg13g2_fill_1 FILLER_63_902 ();
 sg13g2_decap_4 FILLER_63_927 ();
 sg13g2_fill_1 FILLER_63_931 ();
 sg13g2_fill_2 FILLER_63_941 ();
 sg13g2_fill_1 FILLER_63_943 ();
 sg13g2_decap_8 FILLER_63_1013 ();
 sg13g2_decap_8 FILLER_63_1020 ();
 sg13g2_fill_2 FILLER_63_1027 ();
 sg13g2_fill_2 FILLER_64_41 ();
 sg13g2_fill_1 FILLER_64_43 ();
 sg13g2_fill_1 FILLER_64_71 ();
 sg13g2_fill_2 FILLER_64_86 ();
 sg13g2_fill_1 FILLER_64_88 ();
 sg13g2_fill_2 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_130 ();
 sg13g2_decap_4 FILLER_64_137 ();
 sg13g2_fill_1 FILLER_64_141 ();
 sg13g2_fill_1 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_178 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_fill_2 FILLER_64_186 ();
 sg13g2_fill_1 FILLER_64_188 ();
 sg13g2_decap_4 FILLER_64_242 ();
 sg13g2_fill_1 FILLER_64_246 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_4 FILLER_64_313 ();
 sg13g2_fill_2 FILLER_64_326 ();
 sg13g2_decap_8 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_339 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_2 FILLER_64_347 ();
 sg13g2_fill_1 FILLER_64_349 ();
 sg13g2_fill_1 FILLER_64_358 ();
 sg13g2_fill_1 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_429 ();
 sg13g2_decap_8 FILLER_64_459 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_fill_1 FILLER_64_473 ();
 sg13g2_fill_2 FILLER_64_485 ();
 sg13g2_decap_4 FILLER_64_508 ();
 sg13g2_decap_4 FILLER_64_550 ();
 sg13g2_fill_2 FILLER_64_554 ();
 sg13g2_decap_8 FILLER_64_588 ();
 sg13g2_fill_2 FILLER_64_636 ();
 sg13g2_fill_2 FILLER_64_665 ();
 sg13g2_fill_2 FILLER_64_694 ();
 sg13g2_fill_2 FILLER_64_746 ();
 sg13g2_fill_1 FILLER_64_748 ();
 sg13g2_decap_4 FILLER_64_770 ();
 sg13g2_fill_1 FILLER_64_774 ();
 sg13g2_fill_1 FILLER_64_794 ();
 sg13g2_fill_1 FILLER_64_821 ();
 sg13g2_decap_4 FILLER_64_827 ();
 sg13g2_fill_1 FILLER_64_831 ();
 sg13g2_decap_4 FILLER_64_858 ();
 sg13g2_decap_8 FILLER_64_883 ();
 sg13g2_fill_2 FILLER_64_890 ();
 sg13g2_decap_8 FILLER_64_896 ();
 sg13g2_fill_2 FILLER_64_903 ();
 sg13g2_fill_1 FILLER_64_905 ();
 sg13g2_fill_1 FILLER_64_917 ();
 sg13g2_decap_8 FILLER_64_945 ();
 sg13g2_decap_4 FILLER_64_952 ();
 sg13g2_fill_1 FILLER_64_956 ();
 sg13g2_fill_2 FILLER_65_42 ();
 sg13g2_fill_2 FILLER_65_66 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_decap_4 FILLER_65_110 ();
 sg13g2_fill_1 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_4 FILLER_65_140 ();
 sg13g2_fill_2 FILLER_65_144 ();
 sg13g2_decap_4 FILLER_65_164 ();
 sg13g2_decap_4 FILLER_65_172 ();
 sg13g2_fill_2 FILLER_65_176 ();
 sg13g2_fill_2 FILLER_65_183 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_207 ();
 sg13g2_decap_8 FILLER_65_214 ();
 sg13g2_fill_2 FILLER_65_227 ();
 sg13g2_fill_1 FILLER_65_229 ();
 sg13g2_decap_8 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_247 ();
 sg13g2_decap_8 FILLER_65_253 ();
 sg13g2_decap_4 FILLER_65_260 ();
 sg13g2_fill_2 FILLER_65_268 ();
 sg13g2_fill_1 FILLER_65_270 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_353 ();
 sg13g2_decap_4 FILLER_65_359 ();
 sg13g2_decap_8 FILLER_65_377 ();
 sg13g2_decap_8 FILLER_65_384 ();
 sg13g2_fill_2 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_414 ();
 sg13g2_fill_1 FILLER_65_416 ();
 sg13g2_fill_1 FILLER_65_430 ();
 sg13g2_fill_2 FILLER_65_452 ();
 sg13g2_decap_8 FILLER_65_464 ();
 sg13g2_decap_8 FILLER_65_471 ();
 sg13g2_decap_8 FILLER_65_478 ();
 sg13g2_decap_8 FILLER_65_485 ();
 sg13g2_decap_8 FILLER_65_492 ();
 sg13g2_decap_8 FILLER_65_499 ();
 sg13g2_fill_2 FILLER_65_506 ();
 sg13g2_decap_8 FILLER_65_521 ();
 sg13g2_decap_8 FILLER_65_528 ();
 sg13g2_decap_8 FILLER_65_535 ();
 sg13g2_decap_8 FILLER_65_542 ();
 sg13g2_fill_2 FILLER_65_549 ();
 sg13g2_fill_2 FILLER_65_564 ();
 sg13g2_decap_4 FILLER_65_571 ();
 sg13g2_fill_1 FILLER_65_575 ();
 sg13g2_decap_8 FILLER_65_589 ();
 sg13g2_decap_8 FILLER_65_596 ();
 sg13g2_fill_1 FILLER_65_603 ();
 sg13g2_decap_4 FILLER_65_617 ();
 sg13g2_fill_1 FILLER_65_621 ();
 sg13g2_decap_8 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_642 ();
 sg13g2_fill_2 FILLER_65_656 ();
 sg13g2_fill_2 FILLER_65_765 ();
 sg13g2_decap_8 FILLER_65_771 ();
 sg13g2_decap_4 FILLER_65_778 ();
 sg13g2_fill_2 FILLER_65_782 ();
 sg13g2_fill_2 FILLER_65_885 ();
 sg13g2_fill_1 FILLER_65_887 ();
 sg13g2_fill_1 FILLER_65_909 ();
 sg13g2_fill_2 FILLER_65_916 ();
 sg13g2_fill_1 FILLER_65_918 ();
 sg13g2_decap_4 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_955 ();
 sg13g2_decap_8 FILLER_65_962 ();
 sg13g2_decap_4 FILLER_65_969 ();
 sg13g2_fill_1 FILLER_65_973 ();
 sg13g2_decap_4 FILLER_65_1024 ();
 sg13g2_fill_1 FILLER_65_1028 ();
 sg13g2_fill_2 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_2 ();
 sg13g2_fill_1 FILLER_66_30 ();
 sg13g2_fill_2 FILLER_66_45 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_decap_8 FILLER_66_58 ();
 sg13g2_decap_4 FILLER_66_116 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_fill_1 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_186 ();
 sg13g2_fill_1 FILLER_66_188 ();
 sg13g2_decap_8 FILLER_66_193 ();
 sg13g2_decap_4 FILLER_66_200 ();
 sg13g2_fill_2 FILLER_66_204 ();
 sg13g2_decap_8 FILLER_66_221 ();
 sg13g2_decap_4 FILLER_66_228 ();
 sg13g2_fill_2 FILLER_66_232 ();
 sg13g2_fill_2 FILLER_66_252 ();
 sg13g2_fill_2 FILLER_66_264 ();
 sg13g2_fill_2 FILLER_66_283 ();
 sg13g2_fill_1 FILLER_66_285 ();
 sg13g2_fill_2 FILLER_66_295 ();
 sg13g2_fill_1 FILLER_66_297 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_335 ();
 sg13g2_fill_1 FILLER_66_337 ();
 sg13g2_decap_8 FILLER_66_363 ();
 sg13g2_decap_8 FILLER_66_370 ();
 sg13g2_decap_8 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_fill_2 FILLER_66_391 ();
 sg13g2_fill_1 FILLER_66_393 ();
 sg13g2_fill_2 FILLER_66_411 ();
 sg13g2_fill_1 FILLER_66_413 ();
 sg13g2_fill_2 FILLER_66_418 ();
 sg13g2_fill_1 FILLER_66_420 ();
 sg13g2_fill_1 FILLER_66_448 ();
 sg13g2_fill_1 FILLER_66_467 ();
 sg13g2_fill_1 FILLER_66_496 ();
 sg13g2_decap_8 FILLER_66_525 ();
 sg13g2_decap_8 FILLER_66_532 ();
 sg13g2_fill_2 FILLER_66_539 ();
 sg13g2_fill_2 FILLER_66_572 ();
 sg13g2_decap_8 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_fill_1 FILLER_66_602 ();
 sg13g2_decap_4 FILLER_66_631 ();
 sg13g2_fill_1 FILLER_66_689 ();
 sg13g2_fill_1 FILLER_66_733 ();
 sg13g2_decap_8 FILLER_66_761 ();
 sg13g2_decap_8 FILLER_66_768 ();
 sg13g2_fill_1 FILLER_66_775 ();
 sg13g2_fill_2 FILLER_66_781 ();
 sg13g2_fill_1 FILLER_66_783 ();
 sg13g2_decap_8 FILLER_66_816 ();
 sg13g2_decap_4 FILLER_66_836 ();
 sg13g2_fill_2 FILLER_66_840 ();
 sg13g2_fill_2 FILLER_66_869 ();
 sg13g2_fill_2 FILLER_66_879 ();
 sg13g2_decap_4 FILLER_66_886 ();
 sg13g2_fill_2 FILLER_66_890 ();
 sg13g2_fill_1 FILLER_66_913 ();
 sg13g2_decap_4 FILLER_66_950 ();
 sg13g2_fill_1 FILLER_66_954 ();
 sg13g2_fill_2 FILLER_66_966 ();
 sg13g2_fill_1 FILLER_66_968 ();
 sg13g2_decap_4 FILLER_66_988 ();
 sg13g2_decap_4 FILLER_66_1023 ();
 sg13g2_fill_2 FILLER_66_1027 ();
 sg13g2_decap_8 FILLER_67_4 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_65 ();
 sg13g2_decap_4 FILLER_67_72 ();
 sg13g2_fill_2 FILLER_67_76 ();
 sg13g2_fill_2 FILLER_67_107 ();
 sg13g2_fill_2 FILLER_67_128 ();
 sg13g2_fill_1 FILLER_67_166 ();
 sg13g2_fill_2 FILLER_67_193 ();
 sg13g2_fill_1 FILLER_67_195 ();
 sg13g2_decap_8 FILLER_67_228 ();
 sg13g2_decap_4 FILLER_67_235 ();
 sg13g2_fill_1 FILLER_67_239 ();
 sg13g2_fill_2 FILLER_67_252 ();
 sg13g2_fill_1 FILLER_67_254 ();
 sg13g2_fill_1 FILLER_67_260 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_268 ();
 sg13g2_fill_2 FILLER_67_275 ();
 sg13g2_fill_2 FILLER_67_318 ();
 sg13g2_fill_1 FILLER_67_320 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_fill_1 FILLER_67_409 ();
 sg13g2_decap_4 FILLER_67_416 ();
 sg13g2_fill_2 FILLER_67_420 ();
 sg13g2_fill_2 FILLER_67_437 ();
 sg13g2_fill_2 FILLER_67_478 ();
 sg13g2_decap_4 FILLER_67_489 ();
 sg13g2_fill_2 FILLER_67_493 ();
 sg13g2_fill_2 FILLER_67_504 ();
 sg13g2_fill_1 FILLER_67_506 ();
 sg13g2_fill_1 FILLER_67_520 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_fill_1 FILLER_67_589 ();
 sg13g2_fill_2 FILLER_67_621 ();
 sg13g2_fill_1 FILLER_67_690 ();
 sg13g2_fill_2 FILLER_67_747 ();
 sg13g2_fill_1 FILLER_67_749 ();
 sg13g2_fill_2 FILLER_67_769 ();
 sg13g2_fill_1 FILLER_67_771 ();
 sg13g2_fill_2 FILLER_67_800 ();
 sg13g2_fill_2 FILLER_67_839 ();
 sg13g2_fill_1 FILLER_67_841 ();
 sg13g2_decap_8 FILLER_67_848 ();
 sg13g2_decap_4 FILLER_67_855 ();
 sg13g2_fill_1 FILLER_67_859 ();
 sg13g2_fill_2 FILLER_67_869 ();
 sg13g2_fill_1 FILLER_67_871 ();
 sg13g2_fill_2 FILLER_67_884 ();
 sg13g2_decap_8 FILLER_67_908 ();
 sg13g2_fill_1 FILLER_67_915 ();
 sg13g2_fill_1 FILLER_67_943 ();
 sg13g2_decap_8 FILLER_67_957 ();
 sg13g2_decap_8 FILLER_67_964 ();
 sg13g2_decap_4 FILLER_67_971 ();
 sg13g2_fill_1 FILLER_67_1028 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_28 ();
 sg13g2_fill_1 FILLER_68_30 ();
 sg13g2_fill_1 FILLER_68_40 ();
 sg13g2_decap_4 FILLER_68_140 ();
 sg13g2_fill_2 FILLER_68_144 ();
 sg13g2_fill_1 FILLER_68_168 ();
 sg13g2_fill_2 FILLER_68_179 ();
 sg13g2_fill_1 FILLER_68_195 ();
 sg13g2_decap_8 FILLER_68_221 ();
 sg13g2_fill_2 FILLER_68_228 ();
 sg13g2_fill_2 FILLER_68_298 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_fill_2 FILLER_68_321 ();
 sg13g2_fill_1 FILLER_68_323 ();
 sg13g2_fill_1 FILLER_68_337 ();
 sg13g2_decap_8 FILLER_68_342 ();
 sg13g2_decap_4 FILLER_68_349 ();
 sg13g2_decap_8 FILLER_68_361 ();
 sg13g2_fill_2 FILLER_68_368 ();
 sg13g2_fill_1 FILLER_68_370 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_2 FILLER_68_395 ();
 sg13g2_fill_1 FILLER_68_397 ();
 sg13g2_fill_2 FILLER_68_411 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_fill_1 FILLER_68_430 ();
 sg13g2_decap_4 FILLER_68_452 ();
 sg13g2_fill_2 FILLER_68_464 ();
 sg13g2_fill_1 FILLER_68_466 ();
 sg13g2_fill_2 FILLER_68_479 ();
 sg13g2_fill_1 FILLER_68_481 ();
 sg13g2_fill_2 FILLER_68_496 ();
 sg13g2_fill_2 FILLER_68_548 ();
 sg13g2_fill_2 FILLER_68_562 ();
 sg13g2_fill_1 FILLER_68_564 ();
 sg13g2_fill_1 FILLER_68_585 ();
 sg13g2_decap_8 FILLER_68_604 ();
 sg13g2_decap_8 FILLER_68_628 ();
 sg13g2_decap_8 FILLER_68_657 ();
 sg13g2_decap_4 FILLER_68_664 ();
 sg13g2_decap_8 FILLER_68_673 ();
 sg13g2_decap_8 FILLER_68_680 ();
 sg13g2_decap_8 FILLER_68_687 ();
 sg13g2_fill_1 FILLER_68_694 ();
 sg13g2_decap_8 FILLER_68_708 ();
 sg13g2_decap_4 FILLER_68_715 ();
 sg13g2_fill_2 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_4 FILLER_68_770 ();
 sg13g2_fill_2 FILLER_68_774 ();
 sg13g2_fill_1 FILLER_68_814 ();
 sg13g2_fill_1 FILLER_68_820 ();
 sg13g2_fill_2 FILLER_68_870 ();
 sg13g2_fill_1 FILLER_68_885 ();
 sg13g2_fill_2 FILLER_68_891 ();
 sg13g2_fill_1 FILLER_68_893 ();
 sg13g2_fill_1 FILLER_68_917 ();
 sg13g2_decap_8 FILLER_68_928 ();
 sg13g2_decap_8 FILLER_68_935 ();
 sg13g2_decap_4 FILLER_68_942 ();
 sg13g2_fill_1 FILLER_68_946 ();
 sg13g2_fill_2 FILLER_68_965 ();
 sg13g2_fill_2 FILLER_68_987 ();
 sg13g2_fill_1 FILLER_68_989 ();
 sg13g2_decap_8 FILLER_68_1017 ();
 sg13g2_decap_4 FILLER_68_1024 ();
 sg13g2_fill_1 FILLER_68_1028 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_7 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_39 ();
 sg13g2_fill_1 FILLER_69_41 ();
 sg13g2_fill_2 FILLER_69_61 ();
 sg13g2_decap_4 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_decap_8 FILLER_69_219 ();
 sg13g2_fill_2 FILLER_69_226 ();
 sg13g2_fill_2 FILLER_69_282 ();
 sg13g2_decap_4 FILLER_69_316 ();
 sg13g2_fill_2 FILLER_69_320 ();
 sg13g2_fill_2 FILLER_69_358 ();
 sg13g2_fill_1 FILLER_69_360 ();
 sg13g2_fill_2 FILLER_69_389 ();
 sg13g2_fill_2 FILLER_69_414 ();
 sg13g2_fill_1 FILLER_69_437 ();
 sg13g2_decap_4 FILLER_69_453 ();
 sg13g2_fill_1 FILLER_69_457 ();
 sg13g2_fill_1 FILLER_69_464 ();
 sg13g2_fill_1 FILLER_69_491 ();
 sg13g2_fill_1 FILLER_69_505 ();
 sg13g2_decap_8 FILLER_69_525 ();
 sg13g2_fill_2 FILLER_69_532 ();
 sg13g2_decap_8 FILLER_69_547 ();
 sg13g2_fill_2 FILLER_69_554 ();
 sg13g2_decap_4 FILLER_69_572 ();
 sg13g2_fill_2 FILLER_69_614 ();
 sg13g2_fill_2 FILLER_69_624 ();
 sg13g2_fill_1 FILLER_69_626 ();
 sg13g2_decap_8 FILLER_69_652 ();
 sg13g2_fill_2 FILLER_69_659 ();
 sg13g2_decap_4 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_695 ();
 sg13g2_decap_4 FILLER_69_706 ();
 sg13g2_fill_2 FILLER_69_710 ();
 sg13g2_decap_8 FILLER_69_717 ();
 sg13g2_fill_2 FILLER_69_737 ();
 sg13g2_fill_1 FILLER_69_739 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_decap_4 FILLER_69_756 ();
 sg13g2_fill_1 FILLER_69_760 ();
 sg13g2_decap_8 FILLER_69_774 ();
 sg13g2_fill_2 FILLER_69_789 ();
 sg13g2_fill_1 FILLER_69_791 ();
 sg13g2_decap_4 FILLER_69_805 ();
 sg13g2_fill_2 FILLER_69_809 ();
 sg13g2_fill_1 FILLER_69_870 ();
 sg13g2_fill_1 FILLER_69_894 ();
 sg13g2_fill_1 FILLER_69_913 ();
 sg13g2_fill_2 FILLER_69_920 ();
 sg13g2_fill_1 FILLER_69_922 ();
 sg13g2_fill_2 FILLER_69_962 ();
 sg13g2_decap_8 FILLER_69_995 ();
 sg13g2_decap_4 FILLER_70_4 ();
 sg13g2_fill_2 FILLER_70_22 ();
 sg13g2_fill_1 FILLER_70_39 ();
 sg13g2_fill_1 FILLER_70_60 ();
 sg13g2_decap_4 FILLER_70_104 ();
 sg13g2_decap_4 FILLER_70_150 ();
 sg13g2_fill_1 FILLER_70_154 ();
 sg13g2_decap_4 FILLER_70_230 ();
 sg13g2_fill_2 FILLER_70_243 ();
 sg13g2_fill_1 FILLER_70_245 ();
 sg13g2_fill_2 FILLER_70_291 ();
 sg13g2_decap_8 FILLER_70_314 ();
 sg13g2_fill_2 FILLER_70_321 ();
 sg13g2_fill_1 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_351 ();
 sg13g2_fill_2 FILLER_70_358 ();
 sg13g2_fill_2 FILLER_70_388 ();
 sg13g2_decap_4 FILLER_70_417 ();
 sg13g2_fill_2 FILLER_70_421 ();
 sg13g2_fill_2 FILLER_70_449 ();
 sg13g2_fill_1 FILLER_70_451 ();
 sg13g2_fill_1 FILLER_70_462 ();
 sg13g2_fill_2 FILLER_70_472 ();
 sg13g2_fill_2 FILLER_70_500 ();
 sg13g2_decap_8 FILLER_70_521 ();
 sg13g2_decap_8 FILLER_70_528 ();
 sg13g2_decap_8 FILLER_70_535 ();
 sg13g2_decap_4 FILLER_70_542 ();
 sg13g2_fill_1 FILLER_70_546 ();
 sg13g2_fill_2 FILLER_70_602 ();
 sg13g2_fill_1 FILLER_70_640 ();
 sg13g2_fill_2 FILLER_70_737 ();
 sg13g2_fill_2 FILLER_70_744 ();
 sg13g2_fill_1 FILLER_70_746 ();
 sg13g2_decap_8 FILLER_70_775 ();
 sg13g2_fill_2 FILLER_70_782 ();
 sg13g2_fill_1 FILLER_70_784 ();
 sg13g2_fill_2 FILLER_70_790 ();
 sg13g2_fill_1 FILLER_70_792 ();
 sg13g2_decap_8 FILLER_70_806 ();
 sg13g2_fill_2 FILLER_70_813 ();
 sg13g2_fill_1 FILLER_70_815 ();
 sg13g2_decap_8 FILLER_70_829 ();
 sg13g2_decap_4 FILLER_70_836 ();
 sg13g2_fill_2 FILLER_70_840 ();
 sg13g2_decap_4 FILLER_70_847 ();
 sg13g2_fill_1 FILLER_70_851 ();
 sg13g2_fill_2 FILLER_70_872 ();
 sg13g2_decap_4 FILLER_70_893 ();
 sg13g2_fill_1 FILLER_70_919 ();
 sg13g2_fill_2 FILLER_70_971 ();
 sg13g2_fill_1 FILLER_70_973 ();
 sg13g2_fill_2 FILLER_70_980 ();
 sg13g2_decap_8 FILLER_70_1018 ();
 sg13g2_decap_4 FILLER_70_1025 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_61 ();
 sg13g2_fill_1 FILLER_71_78 ();
 sg13g2_decap_8 FILLER_71_151 ();
 sg13g2_fill_1 FILLER_71_190 ();
 sg13g2_decap_8 FILLER_71_200 ();
 sg13g2_decap_4 FILLER_71_244 ();
 sg13g2_fill_2 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_255 ();
 sg13g2_fill_2 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_324 ();
 sg13g2_decap_8 FILLER_71_334 ();
 sg13g2_decap_4 FILLER_71_341 ();
 sg13g2_fill_2 FILLER_71_345 ();
 sg13g2_fill_2 FILLER_71_360 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_fill_2 FILLER_71_382 ();
 sg13g2_fill_1 FILLER_71_410 ();
 sg13g2_fill_2 FILLER_71_416 ();
 sg13g2_fill_1 FILLER_71_418 ();
 sg13g2_decap_4 FILLER_71_423 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_2 FILLER_71_434 ();
 sg13g2_decap_8 FILLER_71_444 ();
 sg13g2_fill_1 FILLER_71_451 ();
 sg13g2_decap_8 FILLER_71_472 ();
 sg13g2_decap_8 FILLER_71_479 ();
 sg13g2_decap_4 FILLER_71_486 ();
 sg13g2_fill_2 FILLER_71_490 ();
 sg13g2_fill_2 FILLER_71_549 ();
 sg13g2_fill_1 FILLER_71_569 ();
 sg13g2_decap_8 FILLER_71_600 ();
 sg13g2_fill_1 FILLER_71_607 ();
 sg13g2_decap_4 FILLER_71_646 ();
 sg13g2_fill_2 FILLER_71_650 ();
 sg13g2_decap_8 FILLER_71_675 ();
 sg13g2_fill_2 FILLER_71_682 ();
 sg13g2_fill_1 FILLER_71_684 ();
 sg13g2_decap_8 FILLER_71_707 ();
 sg13g2_decap_4 FILLER_71_714 ();
 sg13g2_fill_2 FILLER_71_718 ();
 sg13g2_fill_2 FILLER_71_725 ();
 sg13g2_decap_8 FILLER_71_732 ();
 sg13g2_decap_4 FILLER_71_739 ();
 sg13g2_fill_1 FILLER_71_743 ();
 sg13g2_fill_2 FILLER_71_749 ();
 sg13g2_fill_1 FILLER_71_751 ();
 sg13g2_fill_2 FILLER_71_767 ();
 sg13g2_fill_1 FILLER_71_769 ();
 sg13g2_fill_2 FILLER_71_778 ();
 sg13g2_fill_1 FILLER_71_780 ();
 sg13g2_decap_8 FILLER_71_800 ();
 sg13g2_fill_2 FILLER_71_807 ();
 sg13g2_fill_1 FILLER_71_809 ();
 sg13g2_decap_4 FILLER_71_843 ();
 sg13g2_decap_4 FILLER_71_874 ();
 sg13g2_decap_8 FILLER_71_962 ();
 sg13g2_decap_4 FILLER_71_997 ();
 sg13g2_fill_1 FILLER_71_1028 ();
 sg13g2_decap_8 FILLER_72_59 ();
 sg13g2_fill_1 FILLER_72_66 ();
 sg13g2_fill_2 FILLER_72_174 ();
 sg13g2_fill_1 FILLER_72_176 ();
 sg13g2_decap_8 FILLER_72_186 ();
 sg13g2_decap_8 FILLER_72_193 ();
 sg13g2_decap_8 FILLER_72_200 ();
 sg13g2_decap_8 FILLER_72_220 ();
 sg13g2_decap_8 FILLER_72_227 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_299 ();
 sg13g2_decap_8 FILLER_72_328 ();
 sg13g2_decap_4 FILLER_72_335 ();
 sg13g2_fill_2 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_360 ();
 sg13g2_decap_8 FILLER_72_374 ();
 sg13g2_decap_8 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_388 ();
 sg13g2_fill_1 FILLER_72_390 ();
 sg13g2_fill_2 FILLER_72_437 ();
 sg13g2_fill_1 FILLER_72_439 ();
 sg13g2_fill_1 FILLER_72_453 ();
 sg13g2_decap_4 FILLER_72_471 ();
 sg13g2_fill_2 FILLER_72_483 ();
 sg13g2_decap_8 FILLER_72_495 ();
 sg13g2_decap_4 FILLER_72_502 ();
 sg13g2_fill_1 FILLER_72_506 ();
 sg13g2_decap_4 FILLER_72_520 ();
 sg13g2_fill_2 FILLER_72_541 ();
 sg13g2_fill_1 FILLER_72_570 ();
 sg13g2_fill_2 FILLER_72_580 ();
 sg13g2_decap_8 FILLER_72_590 ();
 sg13g2_decap_4 FILLER_72_597 ();
 sg13g2_fill_1 FILLER_72_601 ();
 sg13g2_fill_1 FILLER_72_618 ();
 sg13g2_fill_2 FILLER_72_635 ();
 sg13g2_decap_8 FILLER_72_646 ();
 sg13g2_fill_2 FILLER_72_653 ();
 sg13g2_fill_1 FILLER_72_660 ();
 sg13g2_decap_8 FILLER_72_677 ();
 sg13g2_fill_2 FILLER_72_684 ();
 sg13g2_fill_1 FILLER_72_686 ();
 sg13g2_fill_1 FILLER_72_698 ();
 sg13g2_fill_1 FILLER_72_708 ();
 sg13g2_fill_2 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_771 ();
 sg13g2_decap_8 FILLER_72_778 ();
 sg13g2_fill_1 FILLER_72_788 ();
 sg13g2_decap_4 FILLER_72_794 ();
 sg13g2_fill_1 FILLER_72_798 ();
 sg13g2_fill_2 FILLER_72_946 ();
 sg13g2_fill_1 FILLER_72_974 ();
 sg13g2_fill_2 FILLER_72_985 ();
 sg13g2_fill_2 FILLER_72_1000 ();
 sg13g2_fill_1 FILLER_72_1002 ();
 sg13g2_decap_8 FILLER_72_1012 ();
 sg13g2_decap_8 FILLER_72_1019 ();
 sg13g2_fill_2 FILLER_72_1026 ();
 sg13g2_fill_1 FILLER_72_1028 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_25 ();
 sg13g2_decap_4 FILLER_73_46 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_fill_2 FILLER_73_102 ();
 sg13g2_fill_2 FILLER_73_137 ();
 sg13g2_decap_8 FILLER_73_157 ();
 sg13g2_fill_1 FILLER_73_164 ();
 sg13g2_decap_4 FILLER_73_211 ();
 sg13g2_fill_1 FILLER_73_215 ();
 sg13g2_fill_2 FILLER_73_278 ();
 sg13g2_fill_1 FILLER_73_280 ();
 sg13g2_decap_4 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_311 ();
 sg13g2_fill_2 FILLER_73_360 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_fill_2 FILLER_73_426 ();
 sg13g2_fill_1 FILLER_73_428 ();
 sg13g2_fill_2 FILLER_73_449 ();
 sg13g2_decap_4 FILLER_73_472 ();
 sg13g2_fill_1 FILLER_73_481 ();
 sg13g2_decap_8 FILLER_73_491 ();
 sg13g2_decap_4 FILLER_73_498 ();
 sg13g2_fill_2 FILLER_73_502 ();
 sg13g2_fill_1 FILLER_73_520 ();
 sg13g2_fill_2 FILLER_73_532 ();
 sg13g2_fill_1 FILLER_73_534 ();
 sg13g2_fill_2 FILLER_73_552 ();
 sg13g2_fill_1 FILLER_73_554 ();
 sg13g2_fill_1 FILLER_73_560 ();
 sg13g2_fill_2 FILLER_73_571 ();
 sg13g2_fill_1 FILLER_73_573 ();
 sg13g2_fill_2 FILLER_73_580 ();
 sg13g2_fill_1 FILLER_73_598 ();
 sg13g2_decap_8 FILLER_73_604 ();
 sg13g2_fill_1 FILLER_73_617 ();
 sg13g2_fill_2 FILLER_73_651 ();
 sg13g2_decap_8 FILLER_73_670 ();
 sg13g2_fill_1 FILLER_73_677 ();
 sg13g2_decap_4 FILLER_73_718 ();
 sg13g2_fill_2 FILLER_73_722 ();
 sg13g2_decap_8 FILLER_73_758 ();
 sg13g2_decap_8 FILLER_73_765 ();
 sg13g2_decap_8 FILLER_73_824 ();
 sg13g2_fill_2 FILLER_73_888 ();
 sg13g2_fill_1 FILLER_73_895 ();
 sg13g2_decap_8 FILLER_73_919 ();
 sg13g2_decap_8 FILLER_73_926 ();
 sg13g2_decap_8 FILLER_73_933 ();
 sg13g2_decap_8 FILLER_73_940 ();
 sg13g2_decap_8 FILLER_73_947 ();
 sg13g2_fill_1 FILLER_73_987 ();
 sg13g2_decap_8 FILLER_73_1015 ();
 sg13g2_decap_8 FILLER_73_1022 ();
 sg13g2_fill_2 FILLER_74_37 ();
 sg13g2_fill_2 FILLER_74_55 ();
 sg13g2_fill_1 FILLER_74_96 ();
 sg13g2_fill_2 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_216 ();
 sg13g2_decap_8 FILLER_74_230 ();
 sg13g2_fill_2 FILLER_74_237 ();
 sg13g2_fill_1 FILLER_74_239 ();
 sg13g2_fill_1 FILLER_74_245 ();
 sg13g2_decap_4 FILLER_74_256 ();
 sg13g2_fill_2 FILLER_74_309 ();
 sg13g2_fill_1 FILLER_74_311 ();
 sg13g2_decap_8 FILLER_74_339 ();
 sg13g2_decap_4 FILLER_74_346 ();
 sg13g2_fill_2 FILLER_74_350 ();
 sg13g2_fill_2 FILLER_74_373 ();
 sg13g2_fill_1 FILLER_74_375 ();
 sg13g2_fill_2 FILLER_74_411 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_decap_4 FILLER_74_422 ();
 sg13g2_decap_4 FILLER_74_439 ();
 sg13g2_fill_2 FILLER_74_443 ();
 sg13g2_fill_2 FILLER_74_462 ();
 sg13g2_fill_2 FILLER_74_469 ();
 sg13g2_fill_1 FILLER_74_471 ();
 sg13g2_fill_2 FILLER_74_478 ();
 sg13g2_fill_1 FILLER_74_480 ();
 sg13g2_decap_8 FILLER_74_491 ();
 sg13g2_decap_4 FILLER_74_498 ();
 sg13g2_fill_1 FILLER_74_520 ();
 sg13g2_fill_1 FILLER_74_529 ();
 sg13g2_decap_4 FILLER_74_547 ();
 sg13g2_fill_1 FILLER_74_563 ();
 sg13g2_fill_1 FILLER_74_579 ();
 sg13g2_decap_8 FILLER_74_588 ();
 sg13g2_decap_8 FILLER_74_595 ();
 sg13g2_decap_4 FILLER_74_602 ();
 sg13g2_decap_4 FILLER_74_615 ();
 sg13g2_decap_8 FILLER_74_627 ();
 sg13g2_decap_8 FILLER_74_634 ();
 sg13g2_decap_4 FILLER_74_641 ();
 sg13g2_fill_1 FILLER_74_661 ();
 sg13g2_fill_2 FILLER_74_670 ();
 sg13g2_fill_1 FILLER_74_672 ();
 sg13g2_decap_4 FILLER_74_681 ();
 sg13g2_decap_4 FILLER_74_697 ();
 sg13g2_decap_8 FILLER_74_706 ();
 sg13g2_decap_8 FILLER_74_713 ();
 sg13g2_decap_8 FILLER_74_720 ();
 sg13g2_decap_8 FILLER_74_727 ();
 sg13g2_fill_2 FILLER_74_734 ();
 sg13g2_decap_8 FILLER_74_753 ();
 sg13g2_decap_8 FILLER_74_760 ();
 sg13g2_fill_1 FILLER_74_767 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_814 ();
 sg13g2_decap_8 FILLER_74_821 ();
 sg13g2_decap_8 FILLER_74_828 ();
 sg13g2_fill_1 FILLER_74_835 ();
 sg13g2_fill_2 FILLER_74_841 ();
 sg13g2_fill_1 FILLER_74_843 ();
 sg13g2_fill_2 FILLER_74_850 ();
 sg13g2_fill_1 FILLER_74_852 ();
 sg13g2_decap_4 FILLER_74_862 ();
 sg13g2_decap_4 FILLER_74_887 ();
 sg13g2_fill_2 FILLER_74_901 ();
 sg13g2_fill_1 FILLER_74_903 ();
 sg13g2_fill_2 FILLER_74_916 ();
 sg13g2_fill_1 FILLER_74_918 ();
 sg13g2_fill_2 FILLER_74_940 ();
 sg13g2_decap_4 FILLER_74_955 ();
 sg13g2_fill_2 FILLER_74_984 ();
 sg13g2_decap_8 FILLER_74_1013 ();
 sg13g2_decap_8 FILLER_74_1020 ();
 sg13g2_fill_2 FILLER_74_1027 ();
 sg13g2_fill_2 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_2 ();
 sg13g2_fill_2 FILLER_75_71 ();
 sg13g2_fill_2 FILLER_75_110 ();
 sg13g2_fill_2 FILLER_75_199 ();
 sg13g2_fill_1 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_239 ();
 sg13g2_fill_1 FILLER_75_246 ();
 sg13g2_decap_4 FILLER_75_274 ();
 sg13g2_fill_2 FILLER_75_289 ();
 sg13g2_decap_4 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_360 ();
 sg13g2_fill_2 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_388 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_fill_2 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_418 ();
 sg13g2_fill_2 FILLER_75_450 ();
 sg13g2_decap_8 FILLER_75_464 ();
 sg13g2_fill_1 FILLER_75_475 ();
 sg13g2_decap_8 FILLER_75_500 ();
 sg13g2_fill_1 FILLER_75_507 ();
 sg13g2_decap_8 FILLER_75_516 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_530 ();
 sg13g2_fill_1 FILLER_75_537 ();
 sg13g2_decap_4 FILLER_75_546 ();
 sg13g2_fill_1 FILLER_75_550 ();
 sg13g2_fill_2 FILLER_75_559 ();
 sg13g2_fill_1 FILLER_75_561 ();
 sg13g2_decap_8 FILLER_75_572 ();
 sg13g2_decap_4 FILLER_75_579 ();
 sg13g2_fill_2 FILLER_75_592 ();
 sg13g2_fill_1 FILLER_75_594 ();
 sg13g2_fill_2 FILLER_75_613 ();
 sg13g2_decap_8 FILLER_75_628 ();
 sg13g2_fill_2 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_675 ();
 sg13g2_fill_2 FILLER_75_682 ();
 sg13g2_fill_1 FILLER_75_684 ();
 sg13g2_decap_4 FILLER_75_688 ();
 sg13g2_fill_2 FILLER_75_692 ();
 sg13g2_decap_8 FILLER_75_706 ();
 sg13g2_decap_8 FILLER_75_713 ();
 sg13g2_decap_4 FILLER_75_720 ();
 sg13g2_fill_2 FILLER_75_724 ();
 sg13g2_fill_2 FILLER_75_743 ();
 sg13g2_decap_4 FILLER_75_758 ();
 sg13g2_fill_1 FILLER_75_762 ();
 sg13g2_decap_4 FILLER_75_767 ();
 sg13g2_fill_1 FILLER_75_771 ();
 sg13g2_fill_2 FILLER_75_787 ();
 sg13g2_decap_4 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_815 ();
 sg13g2_fill_1 FILLER_75_822 ();
 sg13g2_fill_1 FILLER_75_849 ();
 sg13g2_fill_2 FILLER_75_862 ();
 sg13g2_fill_1 FILLER_75_864 ();
 sg13g2_fill_2 FILLER_75_871 ();
 sg13g2_fill_1 FILLER_75_873 ();
 sg13g2_decap_8 FILLER_75_885 ();
 sg13g2_decap_8 FILLER_75_892 ();
 sg13g2_fill_2 FILLER_75_899 ();
 sg13g2_fill_1 FILLER_75_901 ();
 sg13g2_decap_4 FILLER_75_907 ();
 sg13g2_decap_4 FILLER_75_937 ();
 sg13g2_fill_1 FILLER_75_941 ();
 sg13g2_fill_1 FILLER_75_984 ();
 sg13g2_fill_2 FILLER_75_994 ();
 sg13g2_fill_1 FILLER_75_996 ();
 sg13g2_decap_8 FILLER_75_1006 ();
 sg13g2_decap_8 FILLER_75_1013 ();
 sg13g2_decap_8 FILLER_75_1020 ();
 sg13g2_fill_2 FILLER_75_1027 ();
 sg13g2_fill_1 FILLER_76_4 ();
 sg13g2_fill_1 FILLER_76_40 ();
 sg13g2_fill_2 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_109 ();
 sg13g2_fill_2 FILLER_76_122 ();
 sg13g2_fill_2 FILLER_76_136 ();
 sg13g2_fill_1 FILLER_76_138 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_fill_1 FILLER_76_168 ();
 sg13g2_fill_2 FILLER_76_179 ();
 sg13g2_fill_1 FILLER_76_181 ();
 sg13g2_decap_4 FILLER_76_186 ();
 sg13g2_decap_4 FILLER_76_199 ();
 sg13g2_fill_2 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_214 ();
 sg13g2_fill_1 FILLER_76_221 ();
 sg13g2_fill_2 FILLER_76_292 ();
 sg13g2_fill_2 FILLER_76_312 ();
 sg13g2_fill_1 FILLER_76_314 ();
 sg13g2_decap_8 FILLER_76_326 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_decap_4 FILLER_76_375 ();
 sg13g2_fill_2 FILLER_76_379 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_fill_2 FILLER_76_397 ();
 sg13g2_fill_1 FILLER_76_399 ();
 sg13g2_fill_1 FILLER_76_414 ();
 sg13g2_fill_2 FILLER_76_425 ();
 sg13g2_decap_4 FILLER_76_434 ();
 sg13g2_fill_2 FILLER_76_438 ();
 sg13g2_fill_2 FILLER_76_446 ();
 sg13g2_decap_8 FILLER_76_452 ();
 sg13g2_decap_8 FILLER_76_459 ();
 sg13g2_fill_2 FILLER_76_524 ();
 sg13g2_decap_4 FILLER_76_547 ();
 sg13g2_fill_2 FILLER_76_551 ();
 sg13g2_fill_1 FILLER_76_561 ();
 sg13g2_decap_4 FILLER_76_570 ();
 sg13g2_fill_1 FILLER_76_574 ();
 sg13g2_fill_2 FILLER_76_590 ();
 sg13g2_fill_1 FILLER_76_604 ();
 sg13g2_fill_2 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_fill_1 FILLER_76_634 ();
 sg13g2_fill_2 FILLER_76_662 ();
 sg13g2_fill_1 FILLER_76_664 ();
 sg13g2_fill_2 FILLER_76_673 ();
 sg13g2_fill_1 FILLER_76_675 ();
 sg13g2_fill_1 FILLER_76_684 ();
 sg13g2_fill_2 FILLER_76_695 ();
 sg13g2_fill_1 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_4 FILLER_76_723 ();
 sg13g2_decap_4 FILLER_76_732 ();
 sg13g2_fill_1 FILLER_76_746 ();
 sg13g2_fill_1 FILLER_76_755 ();
 sg13g2_fill_2 FILLER_76_811 ();
 sg13g2_fill_1 FILLER_76_813 ();
 sg13g2_fill_2 FILLER_76_905 ();
 sg13g2_fill_2 FILLER_76_946 ();
 sg13g2_fill_1 FILLER_76_948 ();
 sg13g2_decap_8 FILLER_76_976 ();
 sg13g2_decap_8 FILLER_76_983 ();
 sg13g2_decap_8 FILLER_76_990 ();
 sg13g2_decap_8 FILLER_76_997 ();
 sg13g2_decap_8 FILLER_76_1004 ();
 sg13g2_decap_8 FILLER_76_1011 ();
 sg13g2_decap_8 FILLER_76_1018 ();
 sg13g2_decap_4 FILLER_76_1025 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_7 ();
 sg13g2_fill_1 FILLER_77_114 ();
 sg13g2_fill_2 FILLER_77_167 ();
 sg13g2_decap_4 FILLER_77_182 ();
 sg13g2_decap_4 FILLER_77_205 ();
 sg13g2_fill_2 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_258 ();
 sg13g2_fill_2 FILLER_77_337 ();
 sg13g2_fill_1 FILLER_77_339 ();
 sg13g2_decap_8 FILLER_77_367 ();
 sg13g2_fill_1 FILLER_77_374 ();
 sg13g2_decap_4 FILLER_77_394 ();
 sg13g2_fill_1 FILLER_77_398 ();
 sg13g2_fill_1 FILLER_77_412 ();
 sg13g2_decap_4 FILLER_77_437 ();
 sg13g2_fill_1 FILLER_77_441 ();
 sg13g2_fill_2 FILLER_77_461 ();
 sg13g2_decap_4 FILLER_77_476 ();
 sg13g2_fill_1 FILLER_77_480 ();
 sg13g2_fill_2 FILLER_77_511 ();
 sg13g2_fill_1 FILLER_77_513 ();
 sg13g2_decap_8 FILLER_77_519 ();
 sg13g2_fill_2 FILLER_77_556 ();
 sg13g2_fill_1 FILLER_77_558 ();
 sg13g2_fill_1 FILLER_77_571 ();
 sg13g2_fill_1 FILLER_77_590 ();
 sg13g2_fill_1 FILLER_77_607 ();
 sg13g2_decap_8 FILLER_77_621 ();
 sg13g2_fill_2 FILLER_77_628 ();
 sg13g2_fill_2 FILLER_77_691 ();
 sg13g2_fill_1 FILLER_77_693 ();
 sg13g2_fill_1 FILLER_77_704 ();
 sg13g2_fill_1 FILLER_77_718 ();
 sg13g2_fill_2 FILLER_77_728 ();
 sg13g2_fill_1 FILLER_77_730 ();
 sg13g2_fill_2 FILLER_77_744 ();
 sg13g2_fill_1 FILLER_77_751 ();
 sg13g2_fill_2 FILLER_77_760 ();
 sg13g2_fill_1 FILLER_77_762 ();
 sg13g2_fill_2 FILLER_77_778 ();
 sg13g2_fill_1 FILLER_77_780 ();
 sg13g2_fill_2 FILLER_77_792 ();
 sg13g2_fill_1 FILLER_77_794 ();
 sg13g2_decap_4 FILLER_77_808 ();
 sg13g2_decap_8 FILLER_77_817 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_4 FILLER_77_831 ();
 sg13g2_fill_2 FILLER_77_835 ();
 sg13g2_fill_1 FILLER_77_846 ();
 sg13g2_fill_1 FILLER_77_852 ();
 sg13g2_fill_2 FILLER_77_880 ();
 sg13g2_decap_4 FILLER_77_918 ();
 sg13g2_decap_4 FILLER_77_949 ();
 sg13g2_fill_2 FILLER_77_953 ();
 sg13g2_decap_8 FILLER_77_977 ();
 sg13g2_decap_8 FILLER_77_984 ();
 sg13g2_decap_8 FILLER_77_991 ();
 sg13g2_decap_8 FILLER_77_998 ();
 sg13g2_decap_8 FILLER_77_1005 ();
 sg13g2_decap_8 FILLER_77_1012 ();
 sg13g2_decap_8 FILLER_77_1019 ();
 sg13g2_fill_2 FILLER_77_1026 ();
 sg13g2_fill_1 FILLER_77_1028 ();
 sg13g2_fill_2 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_fill_1 FILLER_78_133 ();
 sg13g2_fill_1 FILLER_78_254 ();
 sg13g2_fill_2 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_311 ();
 sg13g2_decap_8 FILLER_78_330 ();
 sg13g2_decap_8 FILLER_78_337 ();
 sg13g2_decap_4 FILLER_78_344 ();
 sg13g2_decap_8 FILLER_78_367 ();
 sg13g2_decap_8 FILLER_78_388 ();
 sg13g2_decap_8 FILLER_78_395 ();
 sg13g2_fill_2 FILLER_78_402 ();
 sg13g2_decap_8 FILLER_78_418 ();
 sg13g2_fill_1 FILLER_78_425 ();
 sg13g2_decap_8 FILLER_78_435 ();
 sg13g2_fill_2 FILLER_78_468 ();
 sg13g2_fill_1 FILLER_78_470 ();
 sg13g2_fill_2 FILLER_78_476 ();
 sg13g2_decap_4 FILLER_78_490 ();
 sg13g2_fill_1 FILLER_78_494 ();
 sg13g2_fill_2 FILLER_78_503 ();
 sg13g2_decap_8 FILLER_78_519 ();
 sg13g2_decap_4 FILLER_78_534 ();
 sg13g2_fill_1 FILLER_78_538 ();
 sg13g2_fill_2 FILLER_78_548 ();
 sg13g2_fill_1 FILLER_78_550 ();
 sg13g2_fill_2 FILLER_78_606 ();
 sg13g2_fill_1 FILLER_78_608 ();
 sg13g2_decap_8 FILLER_78_614 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_fill_1 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_659 ();
 sg13g2_decap_8 FILLER_78_666 ();
 sg13g2_fill_1 FILLER_78_673 ();
 sg13g2_decap_4 FILLER_78_680 ();
 sg13g2_fill_1 FILLER_78_684 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_fill_2 FILLER_78_703 ();
 sg13g2_fill_1 FILLER_78_710 ();
 sg13g2_fill_2 FILLER_78_731 ();
 sg13g2_fill_2 FILLER_78_748 ();
 sg13g2_decap_4 FILLER_78_758 ();
 sg13g2_fill_1 FILLER_78_762 ();
 sg13g2_fill_1 FILLER_78_766 ();
 sg13g2_fill_2 FILLER_78_783 ();
 sg13g2_fill_1 FILLER_78_785 ();
 sg13g2_fill_1 FILLER_78_795 ();
 sg13g2_decap_4 FILLER_78_800 ();
 sg13g2_fill_2 FILLER_78_810 ();
 sg13g2_fill_1 FILLER_78_827 ();
 sg13g2_decap_8 FILLER_78_856 ();
 sg13g2_decap_4 FILLER_78_863 ();
 sg13g2_fill_2 FILLER_78_867 ();
 sg13g2_decap_8 FILLER_78_896 ();
 sg13g2_fill_2 FILLER_78_903 ();
 sg13g2_fill_1 FILLER_78_905 ();
 sg13g2_decap_8 FILLER_78_938 ();
 sg13g2_decap_8 FILLER_78_945 ();
 sg13g2_decap_8 FILLER_78_952 ();
 sg13g2_decap_8 FILLER_78_959 ();
 sg13g2_decap_8 FILLER_78_966 ();
 sg13g2_decap_8 FILLER_78_973 ();
 sg13g2_decap_8 FILLER_78_980 ();
 sg13g2_decap_8 FILLER_78_987 ();
 sg13g2_decap_8 FILLER_78_994 ();
 sg13g2_decap_8 FILLER_78_1001 ();
 sg13g2_decap_8 FILLER_78_1008 ();
 sg13g2_decap_8 FILLER_78_1015 ();
 sg13g2_decap_8 FILLER_78_1022 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_17 ();
 sg13g2_fill_1 FILLER_79_21 ();
 sg13g2_fill_2 FILLER_79_65 ();
 sg13g2_decap_4 FILLER_79_130 ();
 sg13g2_fill_1 FILLER_79_134 ();
 sg13g2_fill_2 FILLER_79_145 ();
 sg13g2_fill_2 FILLER_79_169 ();
 sg13g2_decap_4 FILLER_79_184 ();
 sg13g2_fill_1 FILLER_79_188 ();
 sg13g2_fill_1 FILLER_79_264 ();
 sg13g2_fill_1 FILLER_79_288 ();
 sg13g2_fill_2 FILLER_79_325 ();
 sg13g2_decap_4 FILLER_79_332 ();
 sg13g2_fill_1 FILLER_79_336 ();
 sg13g2_fill_2 FILLER_79_354 ();
 sg13g2_fill_1 FILLER_79_356 ();
 sg13g2_fill_2 FILLER_79_365 ();
 sg13g2_fill_2 FILLER_79_373 ();
 sg13g2_fill_1 FILLER_79_375 ();
 sg13g2_fill_2 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_4 FILLER_79_430 ();
 sg13g2_fill_2 FILLER_79_461 ();
 sg13g2_fill_1 FILLER_79_486 ();
 sg13g2_decap_4 FILLER_79_500 ();
 sg13g2_decap_8 FILLER_79_512 ();
 sg13g2_decap_4 FILLER_79_519 ();
 sg13g2_fill_1 FILLER_79_523 ();
 sg13g2_decap_8 FILLER_79_552 ();
 sg13g2_fill_1 FILLER_79_559 ();
 sg13g2_decap_4 FILLER_79_564 ();
 sg13g2_fill_2 FILLER_79_591 ();
 sg13g2_fill_1 FILLER_79_625 ();
 sg13g2_decap_8 FILLER_79_633 ();
 sg13g2_fill_2 FILLER_79_650 ();
 sg13g2_decap_8 FILLER_79_656 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_4 FILLER_79_676 ();
 sg13g2_fill_2 FILLER_79_680 ();
 sg13g2_decap_8 FILLER_79_695 ();
 sg13g2_fill_2 FILLER_79_702 ();
 sg13g2_fill_2 FILLER_79_719 ();
 sg13g2_fill_2 FILLER_79_726 ();
 sg13g2_fill_1 FILLER_79_728 ();
 sg13g2_decap_4 FILLER_79_758 ();
 sg13g2_decap_4 FILLER_79_770 ();
 sg13g2_fill_2 FILLER_79_774 ();
 sg13g2_fill_2 FILLER_79_781 ();
 sg13g2_fill_1 FILLER_79_783 ();
 sg13g2_decap_4 FILLER_79_788 ();
 sg13g2_fill_2 FILLER_79_802 ();
 sg13g2_fill_1 FILLER_79_804 ();
 sg13g2_decap_4 FILLER_79_818 ();
 sg13g2_decap_4 FILLER_79_850 ();
 sg13g2_fill_2 FILLER_79_854 ();
 sg13g2_decap_4 FILLER_79_869 ();
 sg13g2_decap_8 FILLER_79_886 ();
 sg13g2_decap_8 FILLER_79_893 ();
 sg13g2_fill_1 FILLER_79_900 ();
 sg13g2_decap_8 FILLER_79_937 ();
 sg13g2_decap_8 FILLER_79_944 ();
 sg13g2_decap_8 FILLER_79_951 ();
 sg13g2_decap_8 FILLER_79_958 ();
 sg13g2_decap_8 FILLER_79_965 ();
 sg13g2_decap_8 FILLER_79_972 ();
 sg13g2_decap_8 FILLER_79_979 ();
 sg13g2_decap_8 FILLER_79_986 ();
 sg13g2_decap_8 FILLER_79_993 ();
 sg13g2_decap_8 FILLER_79_1000 ();
 sg13g2_decap_8 FILLER_79_1007 ();
 sg13g2_decap_8 FILLER_79_1014 ();
 sg13g2_decap_8 FILLER_79_1021 ();
 sg13g2_fill_1 FILLER_79_1028 ();
 sg13g2_decap_4 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_4 ();
 sg13g2_fill_1 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_fill_1 FILLER_80_168 ();
 sg13g2_fill_1 FILLER_80_196 ();
 sg13g2_decap_4 FILLER_80_295 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_fill_1 FILLER_80_327 ();
 sg13g2_decap_4 FILLER_80_336 ();
 sg13g2_fill_2 FILLER_80_351 ();
 sg13g2_fill_1 FILLER_80_353 ();
 sg13g2_fill_2 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_4 FILLER_80_394 ();
 sg13g2_fill_2 FILLER_80_402 ();
 sg13g2_fill_1 FILLER_80_404 ();
 sg13g2_decap_8 FILLER_80_410 ();
 sg13g2_fill_1 FILLER_80_450 ();
 sg13g2_decap_4 FILLER_80_464 ();
 sg13g2_decap_8 FILLER_80_489 ();
 sg13g2_fill_2 FILLER_80_496 ();
 sg13g2_decap_8 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_fill_2 FILLER_80_540 ();
 sg13g2_fill_1 FILLER_80_542 ();
 sg13g2_decap_8 FILLER_80_551 ();
 sg13g2_fill_1 FILLER_80_558 ();
 sg13g2_decap_8 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_580 ();
 sg13g2_decap_8 FILLER_80_587 ();
 sg13g2_fill_2 FILLER_80_622 ();
 sg13g2_fill_2 FILLER_80_635 ();
 sg13g2_fill_2 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_683 ();
 sg13g2_fill_2 FILLER_80_690 ();
 sg13g2_fill_1 FILLER_80_697 ();
 sg13g2_decap_4 FILLER_80_715 ();
 sg13g2_fill_1 FILLER_80_719 ();
 sg13g2_fill_2 FILLER_80_724 ();
 sg13g2_fill_1 FILLER_80_726 ();
 sg13g2_fill_2 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_762 ();
 sg13g2_fill_2 FILLER_80_769 ();
 sg13g2_fill_1 FILLER_80_771 ();
 sg13g2_fill_1 FILLER_80_780 ();
 sg13g2_fill_2 FILLER_80_795 ();
 sg13g2_decap_8 FILLER_80_816 ();
 sg13g2_decap_8 FILLER_80_823 ();
 sg13g2_decap_4 FILLER_80_830 ();
 sg13g2_fill_2 FILLER_80_834 ();
 sg13g2_fill_2 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_81_0 ();
 sg13g2_fill_2 FILLER_81_7 ();
 sg13g2_fill_1 FILLER_81_22 ();
 sg13g2_fill_1 FILLER_81_32 ();
 sg13g2_fill_1 FILLER_81_100 ();
 sg13g2_fill_2 FILLER_81_114 ();
 sg13g2_fill_1 FILLER_81_116 ();
 sg13g2_fill_1 FILLER_81_166 ();
 sg13g2_decap_4 FILLER_81_177 ();
 sg13g2_fill_2 FILLER_81_181 ();
 sg13g2_decap_4 FILLER_81_230 ();
 sg13g2_fill_1 FILLER_81_234 ();
 sg13g2_decap_4 FILLER_81_288 ();
 sg13g2_fill_1 FILLER_81_292 ();
 sg13g2_decap_4 FILLER_81_319 ();
 sg13g2_fill_1 FILLER_81_323 ();
 sg13g2_decap_8 FILLER_81_344 ();
 sg13g2_fill_1 FILLER_81_351 ();
 sg13g2_fill_1 FILLER_81_372 ();
 sg13g2_decap_8 FILLER_81_386 ();
 sg13g2_decap_8 FILLER_81_419 ();
 sg13g2_fill_1 FILLER_81_426 ();
 sg13g2_fill_2 FILLER_81_446 ();
 sg13g2_decap_8 FILLER_81_461 ();
 sg13g2_fill_2 FILLER_81_468 ();
 sg13g2_fill_1 FILLER_81_470 ();
 sg13g2_decap_8 FILLER_81_479 ();
 sg13g2_decap_8 FILLER_81_486 ();
 sg13g2_decap_4 FILLER_81_493 ();
 sg13g2_fill_2 FILLER_81_497 ();
 sg13g2_fill_2 FILLER_81_522 ();
 sg13g2_fill_1 FILLER_81_524 ();
 sg13g2_decap_4 FILLER_81_533 ();
 sg13g2_fill_1 FILLER_81_537 ();
 sg13g2_fill_2 FILLER_81_546 ();
 sg13g2_fill_1 FILLER_81_548 ();
 sg13g2_fill_1 FILLER_81_670 ();
 sg13g2_decap_8 FILLER_81_684 ();
 sg13g2_fill_2 FILLER_81_691 ();
 sg13g2_decap_8 FILLER_81_711 ();
 sg13g2_fill_2 FILLER_81_718 ();
 sg13g2_decap_4 FILLER_81_737 ();
 sg13g2_fill_2 FILLER_81_741 ();
 sg13g2_decap_8 FILLER_81_748 ();
 sg13g2_decap_8 FILLER_81_755 ();
 sg13g2_decap_4 FILLER_81_762 ();
 sg13g2_fill_2 FILLER_81_794 ();
 sg13g2_fill_1 FILLER_81_796 ();
 sg13g2_decap_8 FILLER_81_844 ();
 sg13g2_decap_8 FILLER_81_851 ();
 sg13g2_decap_8 FILLER_81_858 ();
 sg13g2_decap_8 FILLER_81_865 ();
 sg13g2_decap_8 FILLER_81_872 ();
 sg13g2_decap_8 FILLER_81_879 ();
 sg13g2_decap_8 FILLER_81_886 ();
 sg13g2_decap_8 FILLER_81_893 ();
 sg13g2_decap_8 FILLER_81_900 ();
 sg13g2_decap_8 FILLER_81_907 ();
 sg13g2_decap_8 FILLER_81_914 ();
 sg13g2_decap_8 FILLER_81_921 ();
 sg13g2_decap_8 FILLER_81_928 ();
 sg13g2_decap_8 FILLER_81_935 ();
 sg13g2_decap_8 FILLER_81_942 ();
 sg13g2_decap_8 FILLER_81_949 ();
 sg13g2_decap_8 FILLER_81_956 ();
 sg13g2_decap_8 FILLER_81_963 ();
 sg13g2_decap_8 FILLER_81_970 ();
 sg13g2_decap_8 FILLER_81_977 ();
 sg13g2_decap_8 FILLER_81_984 ();
 sg13g2_decap_8 FILLER_81_991 ();
 sg13g2_decap_8 FILLER_81_998 ();
 sg13g2_decap_8 FILLER_81_1005 ();
 sg13g2_decap_8 FILLER_81_1012 ();
 sg13g2_decap_8 FILLER_81_1019 ();
 sg13g2_fill_2 FILLER_81_1026 ();
 sg13g2_fill_1 FILLER_81_1028 ();
 sg13g2_decap_8 FILLER_82_158 ();
 sg13g2_fill_2 FILLER_82_165 ();
 sg13g2_decap_8 FILLER_82_195 ();
 sg13g2_fill_1 FILLER_82_250 ();
 sg13g2_fill_2 FILLER_82_282 ();
 sg13g2_fill_1 FILLER_82_284 ();
 sg13g2_decap_8 FILLER_82_336 ();
 sg13g2_decap_8 FILLER_82_343 ();
 sg13g2_fill_2 FILLER_82_350 ();
 sg13g2_fill_2 FILLER_82_368 ();
 sg13g2_fill_1 FILLER_82_370 ();
 sg13g2_fill_1 FILLER_82_380 ();
 sg13g2_fill_1 FILLER_82_393 ();
 sg13g2_decap_8 FILLER_82_418 ();
 sg13g2_decap_8 FILLER_82_425 ();
 sg13g2_decap_4 FILLER_82_432 ();
 sg13g2_fill_2 FILLER_82_436 ();
 sg13g2_fill_1 FILLER_82_442 ();
 sg13g2_fill_1 FILLER_82_451 ();
 sg13g2_fill_2 FILLER_82_465 ();
 sg13g2_fill_1 FILLER_82_467 ();
 sg13g2_fill_2 FILLER_82_494 ();
 sg13g2_fill_1 FILLER_82_517 ();
 sg13g2_decap_8 FILLER_82_552 ();
 sg13g2_decap_8 FILLER_82_559 ();
 sg13g2_decap_8 FILLER_82_566 ();
 sg13g2_decap_8 FILLER_82_577 ();
 sg13g2_fill_2 FILLER_82_584 ();
 sg13g2_fill_1 FILLER_82_602 ();
 sg13g2_fill_2 FILLER_82_667 ();
 sg13g2_decap_4 FILLER_82_678 ();
 sg13g2_decap_4 FILLER_82_689 ();
 sg13g2_fill_1 FILLER_82_693 ();
 sg13g2_fill_2 FILLER_82_702 ();
 sg13g2_decap_8 FILLER_82_732 ();
 sg13g2_fill_2 FILLER_82_739 ();
 sg13g2_fill_1 FILLER_82_741 ();
 sg13g2_fill_2 FILLER_82_763 ();
 sg13g2_fill_2 FILLER_82_808 ();
 sg13g2_fill_1 FILLER_82_810 ();
 sg13g2_decap_8 FILLER_82_839 ();
 sg13g2_decap_8 FILLER_82_846 ();
 sg13g2_decap_8 FILLER_82_853 ();
 sg13g2_decap_8 FILLER_82_860 ();
 sg13g2_decap_8 FILLER_82_867 ();
 sg13g2_decap_8 FILLER_82_874 ();
 sg13g2_decap_8 FILLER_82_881 ();
 sg13g2_decap_8 FILLER_82_888 ();
 sg13g2_decap_8 FILLER_82_895 ();
 sg13g2_decap_8 FILLER_82_902 ();
 sg13g2_decap_8 FILLER_82_909 ();
 sg13g2_decap_8 FILLER_82_916 ();
 sg13g2_decap_8 FILLER_82_923 ();
 sg13g2_decap_8 FILLER_82_930 ();
 sg13g2_decap_8 FILLER_82_937 ();
 sg13g2_decap_8 FILLER_82_944 ();
 sg13g2_decap_8 FILLER_82_951 ();
 sg13g2_decap_8 FILLER_82_958 ();
 sg13g2_decap_8 FILLER_82_965 ();
 sg13g2_decap_8 FILLER_82_972 ();
 sg13g2_decap_8 FILLER_82_979 ();
 sg13g2_decap_8 FILLER_82_986 ();
 sg13g2_decap_8 FILLER_82_993 ();
 sg13g2_decap_8 FILLER_82_1000 ();
 sg13g2_decap_8 FILLER_82_1007 ();
 sg13g2_decap_8 FILLER_82_1014 ();
 sg13g2_decap_8 FILLER_82_1021 ();
 sg13g2_fill_1 FILLER_82_1028 ();
 sg13g2_decap_4 FILLER_83_0 ();
 sg13g2_fill_2 FILLER_83_4 ();
 sg13g2_fill_2 FILLER_83_19 ();
 sg13g2_decap_4 FILLER_83_30 ();
 sg13g2_fill_1 FILLER_83_34 ();
 sg13g2_fill_2 FILLER_83_62 ();
 sg13g2_fill_1 FILLER_83_73 ();
 sg13g2_decap_4 FILLER_83_158 ();
 sg13g2_decap_8 FILLER_83_199 ();
 sg13g2_fill_1 FILLER_83_206 ();
 sg13g2_decap_8 FILLER_83_234 ();
 sg13g2_fill_1 FILLER_83_260 ();
 sg13g2_decap_8 FILLER_83_275 ();
 sg13g2_fill_1 FILLER_83_282 ();
 sg13g2_fill_2 FILLER_83_296 ();
 sg13g2_fill_2 FILLER_83_307 ();
 sg13g2_fill_1 FILLER_83_309 ();
 sg13g2_decap_8 FILLER_83_327 ();
 sg13g2_fill_2 FILLER_83_334 ();
 sg13g2_decap_8 FILLER_83_387 ();
 sg13g2_decap_4 FILLER_83_394 ();
 sg13g2_decap_4 FILLER_83_433 ();
 sg13g2_decap_4 FILLER_83_442 ();
 sg13g2_fill_1 FILLER_83_446 ();
 sg13g2_fill_2 FILLER_83_455 ();
 sg13g2_fill_2 FILLER_83_465 ();
 sg13g2_decap_8 FILLER_83_518 ();
 sg13g2_decap_8 FILLER_83_525 ();
 sg13g2_fill_2 FILLER_83_532 ();
 sg13g2_decap_8 FILLER_83_542 ();
 sg13g2_decap_8 FILLER_83_549 ();
 sg13g2_fill_2 FILLER_83_556 ();
 sg13g2_decap_8 FILLER_83_565 ();
 sg13g2_decap_8 FILLER_83_580 ();
 sg13g2_decap_8 FILLER_83_587 ();
 sg13g2_decap_8 FILLER_83_594 ();
 sg13g2_fill_1 FILLER_83_601 ();
 sg13g2_decap_8 FILLER_83_608 ();
 sg13g2_decap_8 FILLER_83_615 ();
 sg13g2_decap_8 FILLER_83_622 ();
 sg13g2_decap_8 FILLER_83_629 ();
 sg13g2_decap_8 FILLER_83_636 ();
 sg13g2_decap_8 FILLER_83_643 ();
 sg13g2_decap_4 FILLER_83_650 ();
 sg13g2_fill_2 FILLER_83_654 ();
 sg13g2_fill_2 FILLER_83_664 ();
 sg13g2_decap_4 FILLER_83_679 ();
 sg13g2_fill_1 FILLER_83_683 ();
 sg13g2_decap_8 FILLER_83_692 ();
 sg13g2_decap_8 FILLER_83_699 ();
 sg13g2_fill_1 FILLER_83_706 ();
 sg13g2_fill_2 FILLER_83_729 ();
 sg13g2_fill_1 FILLER_83_731 ();
 sg13g2_decap_8 FILLER_83_744 ();
 sg13g2_decap_8 FILLER_83_751 ();
 sg13g2_decap_8 FILLER_83_758 ();
 sg13g2_fill_2 FILLER_83_765 ();
 sg13g2_fill_2 FILLER_83_786 ();
 sg13g2_fill_1 FILLER_83_788 ();
 sg13g2_decap_8 FILLER_83_793 ();
 sg13g2_decap_8 FILLER_83_800 ();
 sg13g2_fill_1 FILLER_83_807 ();
 sg13g2_decap_8 FILLER_83_814 ();
 sg13g2_decap_8 FILLER_83_821 ();
 sg13g2_fill_2 FILLER_83_828 ();
 sg13g2_fill_1 FILLER_83_830 ();
 sg13g2_decap_8 FILLER_83_844 ();
 sg13g2_decap_8 FILLER_83_851 ();
 sg13g2_decap_8 FILLER_83_858 ();
 sg13g2_decap_8 FILLER_83_865 ();
 sg13g2_decap_8 FILLER_83_872 ();
 sg13g2_decap_8 FILLER_83_879 ();
 sg13g2_decap_8 FILLER_83_886 ();
 sg13g2_decap_8 FILLER_83_893 ();
 sg13g2_decap_8 FILLER_83_900 ();
 sg13g2_decap_8 FILLER_83_907 ();
 sg13g2_decap_8 FILLER_83_914 ();
 sg13g2_decap_8 FILLER_83_921 ();
 sg13g2_decap_8 FILLER_83_928 ();
 sg13g2_decap_8 FILLER_83_935 ();
 sg13g2_decap_8 FILLER_83_942 ();
 sg13g2_decap_8 FILLER_83_949 ();
 sg13g2_decap_8 FILLER_83_956 ();
 sg13g2_decap_8 FILLER_83_963 ();
 sg13g2_decap_8 FILLER_83_970 ();
 sg13g2_decap_8 FILLER_83_977 ();
 sg13g2_decap_8 FILLER_83_984 ();
 sg13g2_decap_8 FILLER_83_991 ();
 sg13g2_decap_8 FILLER_83_998 ();
 sg13g2_decap_8 FILLER_83_1005 ();
 sg13g2_decap_8 FILLER_83_1012 ();
 sg13g2_decap_8 FILLER_83_1019 ();
 sg13g2_fill_2 FILLER_83_1026 ();
 sg13g2_fill_1 FILLER_83_1028 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_fill_2 FILLER_84_7 ();
 sg13g2_fill_1 FILLER_84_9 ();
 sg13g2_decap_8 FILLER_84_27 ();
 sg13g2_decap_8 FILLER_84_34 ();
 sg13g2_fill_1 FILLER_84_203 ();
 sg13g2_fill_1 FILLER_84_226 ();
 sg13g2_decap_8 FILLER_84_249 ();
 sg13g2_fill_2 FILLER_84_256 ();
 sg13g2_fill_1 FILLER_84_273 ();
 sg13g2_decap_8 FILLER_84_287 ();
 sg13g2_decap_4 FILLER_84_300 ();
 sg13g2_decap_8 FILLER_84_323 ();
 sg13g2_decap_8 FILLER_84_356 ();
 sg13g2_fill_1 FILLER_84_363 ();
 sg13g2_fill_1 FILLER_84_390 ();
 sg13g2_fill_2 FILLER_84_399 ();
 sg13g2_decap_4 FILLER_84_448 ();
 sg13g2_fill_2 FILLER_84_452 ();
 sg13g2_decap_8 FILLER_84_463 ();
 sg13g2_decap_4 FILLER_84_470 ();
 sg13g2_fill_2 FILLER_84_474 ();
 sg13g2_decap_8 FILLER_84_494 ();
 sg13g2_fill_2 FILLER_84_501 ();
 sg13g2_fill_1 FILLER_84_506 ();
 sg13g2_fill_2 FILLER_84_528 ();
 sg13g2_fill_1 FILLER_84_530 ();
 sg13g2_decap_8 FILLER_84_539 ();
 sg13g2_decap_4 FILLER_84_546 ();
 sg13g2_fill_2 FILLER_84_550 ();
 sg13g2_decap_4 FILLER_84_585 ();
 sg13g2_fill_2 FILLER_84_589 ();
 sg13g2_fill_1 FILLER_84_597 ();
 sg13g2_decap_8 FILLER_84_602 ();
 sg13g2_decap_4 FILLER_84_609 ();
 sg13g2_decap_8 FILLER_84_617 ();
 sg13g2_decap_8 FILLER_84_624 ();
 sg13g2_fill_1 FILLER_84_631 ();
 sg13g2_decap_4 FILLER_84_637 ();
 sg13g2_fill_1 FILLER_84_641 ();
 sg13g2_fill_1 FILLER_84_647 ();
 sg13g2_fill_2 FILLER_84_661 ();
 sg13g2_decap_8 FILLER_84_683 ();
 sg13g2_decap_8 FILLER_84_690 ();
 sg13g2_decap_8 FILLER_84_697 ();
 sg13g2_decap_8 FILLER_84_710 ();
 sg13g2_decap_8 FILLER_84_717 ();
 sg13g2_decap_8 FILLER_84_728 ();
 sg13g2_decap_8 FILLER_84_735 ();
 sg13g2_decap_8 FILLER_84_742 ();
 sg13g2_decap_4 FILLER_84_749 ();
 sg13g2_fill_1 FILLER_84_753 ();
 sg13g2_decap_4 FILLER_84_759 ();
 sg13g2_fill_2 FILLER_84_763 ();
 sg13g2_fill_1 FILLER_84_792 ();
 sg13g2_decap_8 FILLER_84_801 ();
 sg13g2_fill_1 FILLER_84_808 ();
 sg13g2_fill_2 FILLER_84_819 ();
 sg13g2_fill_1 FILLER_84_821 ();
 sg13g2_decap_8 FILLER_84_835 ();
 sg13g2_decap_8 FILLER_84_842 ();
 sg13g2_decap_8 FILLER_84_849 ();
 sg13g2_decap_8 FILLER_84_856 ();
 sg13g2_decap_8 FILLER_84_863 ();
 sg13g2_decap_8 FILLER_84_870 ();
 sg13g2_decap_8 FILLER_84_877 ();
 sg13g2_decap_8 FILLER_84_884 ();
 sg13g2_decap_8 FILLER_84_891 ();
 sg13g2_decap_8 FILLER_84_898 ();
 sg13g2_decap_8 FILLER_84_905 ();
 sg13g2_decap_8 FILLER_84_912 ();
 sg13g2_decap_8 FILLER_84_919 ();
 sg13g2_decap_8 FILLER_84_926 ();
 sg13g2_decap_8 FILLER_84_933 ();
 sg13g2_decap_8 FILLER_84_940 ();
 sg13g2_decap_8 FILLER_84_947 ();
 sg13g2_decap_8 FILLER_84_954 ();
 sg13g2_decap_8 FILLER_84_961 ();
 sg13g2_decap_8 FILLER_84_968 ();
 sg13g2_decap_8 FILLER_84_975 ();
 sg13g2_decap_8 FILLER_84_982 ();
 sg13g2_decap_8 FILLER_84_989 ();
 sg13g2_decap_8 FILLER_84_996 ();
 sg13g2_decap_8 FILLER_84_1003 ();
 sg13g2_decap_8 FILLER_84_1010 ();
 sg13g2_decap_8 FILLER_84_1017 ();
 sg13g2_decap_4 FILLER_84_1024 ();
 sg13g2_fill_1 FILLER_84_1028 ();
 sg13g2_decap_4 FILLER_85_0 ();
 sg13g2_fill_1 FILLER_85_69 ();
 sg13g2_fill_1 FILLER_85_100 ();
 sg13g2_fill_2 FILLER_85_201 ();
 sg13g2_fill_2 FILLER_85_212 ();
 sg13g2_fill_2 FILLER_85_224 ();
 sg13g2_fill_2 FILLER_85_273 ();
 sg13g2_fill_2 FILLER_85_288 ();
 sg13g2_fill_1 FILLER_85_297 ();
 sg13g2_fill_2 FILLER_85_317 ();
 sg13g2_fill_2 FILLER_85_323 ();
 sg13g2_fill_1 FILLER_85_334 ();
 sg13g2_fill_2 FILLER_85_341 ();
 sg13g2_decap_4 FILLER_85_351 ();
 sg13g2_fill_1 FILLER_85_355 ();
 sg13g2_fill_2 FILLER_85_361 ();
 sg13g2_decap_4 FILLER_85_384 ();
 sg13g2_fill_1 FILLER_85_388 ();
 sg13g2_decap_8 FILLER_85_404 ();
 sg13g2_decap_8 FILLER_85_411 ();
 sg13g2_decap_4 FILLER_85_418 ();
 sg13g2_decap_8 FILLER_85_428 ();
 sg13g2_decap_4 FILLER_85_435 ();
 sg13g2_fill_1 FILLER_85_439 ();
 sg13g2_decap_8 FILLER_85_453 ();
 sg13g2_fill_2 FILLER_85_460 ();
 sg13g2_fill_1 FILLER_85_462 ();
 sg13g2_fill_1 FILLER_85_476 ();
 sg13g2_fill_1 FILLER_85_498 ();
 sg13g2_fill_2 FILLER_85_504 ();
 sg13g2_fill_2 FILLER_85_518 ();
 sg13g2_decap_4 FILLER_85_550 ();
 sg13g2_decap_4 FILLER_85_562 ();
 sg13g2_fill_2 FILLER_85_580 ();
 sg13g2_fill_1 FILLER_85_582 ();
 sg13g2_decap_4 FILLER_85_588 ();
 sg13g2_fill_2 FILLER_85_613 ();
 sg13g2_fill_1 FILLER_85_615 ();
 sg13g2_fill_2 FILLER_85_632 ();
 sg13g2_fill_2 FILLER_85_656 ();
 sg13g2_fill_2 FILLER_85_667 ();
 sg13g2_fill_1 FILLER_85_674 ();
 sg13g2_decap_4 FILLER_85_693 ();
 sg13g2_fill_1 FILLER_85_697 ();
 sg13g2_fill_2 FILLER_85_706 ();
 sg13g2_fill_2 FILLER_85_724 ();
 sg13g2_fill_1 FILLER_85_726 ();
 sg13g2_fill_1 FILLER_85_751 ();
 sg13g2_decap_4 FILLER_85_774 ();
 sg13g2_fill_2 FILLER_85_806 ();
 sg13g2_fill_1 FILLER_85_808 ();
 sg13g2_fill_1 FILLER_85_825 ();
 sg13g2_decap_8 FILLER_85_836 ();
 sg13g2_decap_8 FILLER_85_843 ();
 sg13g2_decap_8 FILLER_85_850 ();
 sg13g2_decap_8 FILLER_85_857 ();
 sg13g2_decap_8 FILLER_85_864 ();
 sg13g2_decap_8 FILLER_85_871 ();
 sg13g2_decap_8 FILLER_85_878 ();
 sg13g2_decap_8 FILLER_85_885 ();
 sg13g2_decap_8 FILLER_85_892 ();
 sg13g2_decap_8 FILLER_85_899 ();
 sg13g2_decap_8 FILLER_85_906 ();
 sg13g2_decap_8 FILLER_85_913 ();
 sg13g2_decap_8 FILLER_85_920 ();
 sg13g2_decap_8 FILLER_85_927 ();
 sg13g2_decap_8 FILLER_85_934 ();
 sg13g2_decap_8 FILLER_85_941 ();
 sg13g2_decap_8 FILLER_85_948 ();
 sg13g2_decap_8 FILLER_85_955 ();
 sg13g2_decap_8 FILLER_85_962 ();
 sg13g2_decap_8 FILLER_85_969 ();
 sg13g2_decap_8 FILLER_85_976 ();
 sg13g2_decap_8 FILLER_85_983 ();
 sg13g2_decap_8 FILLER_85_990 ();
 sg13g2_decap_8 FILLER_85_997 ();
 sg13g2_decap_8 FILLER_85_1004 ();
 sg13g2_decap_8 FILLER_85_1011 ();
 sg13g2_decap_8 FILLER_85_1018 ();
 sg13g2_decap_4 FILLER_85_1025 ();
 sg13g2_decap_8 FILLER_86_0 ();
 sg13g2_fill_1 FILLER_86_7 ();
 sg13g2_decap_8 FILLER_86_29 ();
 sg13g2_fill_2 FILLER_86_36 ();
 sg13g2_decap_8 FILLER_86_47 ();
 sg13g2_fill_2 FILLER_86_54 ();
 sg13g2_fill_2 FILLER_86_59 ();
 sg13g2_fill_2 FILLER_86_105 ();
 sg13g2_fill_2 FILLER_86_137 ();
 sg13g2_fill_1 FILLER_86_167 ();
 sg13g2_decap_4 FILLER_86_205 ();
 sg13g2_fill_2 FILLER_86_209 ();
 sg13g2_fill_2 FILLER_86_231 ();
 sg13g2_decap_8 FILLER_86_273 ();
 sg13g2_fill_2 FILLER_86_280 ();
 sg13g2_decap_8 FILLER_86_313 ();
 sg13g2_decap_8 FILLER_86_320 ();
 sg13g2_decap_4 FILLER_86_327 ();
 sg13g2_fill_2 FILLER_86_331 ();
 sg13g2_decap_8 FILLER_86_353 ();
 sg13g2_decap_8 FILLER_86_360 ();
 sg13g2_fill_2 FILLER_86_367 ();
 sg13g2_fill_1 FILLER_86_378 ();
 sg13g2_fill_2 FILLER_86_385 ();
 sg13g2_decap_8 FILLER_86_410 ();
 sg13g2_fill_2 FILLER_86_417 ();
 sg13g2_decap_8 FILLER_86_429 ();
 sg13g2_fill_2 FILLER_86_436 ();
 sg13g2_fill_2 FILLER_86_454 ();
 sg13g2_decap_4 FILLER_86_488 ();
 sg13g2_fill_2 FILLER_86_500 ();
 sg13g2_fill_1 FILLER_86_502 ();
 sg13g2_fill_1 FILLER_86_511 ();
 sg13g2_fill_2 FILLER_86_525 ();
 sg13g2_fill_1 FILLER_86_556 ();
 sg13g2_fill_2 FILLER_86_569 ();
 sg13g2_fill_1 FILLER_86_571 ();
 sg13g2_fill_1 FILLER_86_588 ();
 sg13g2_decap_8 FILLER_86_617 ();
 sg13g2_decap_8 FILLER_86_624 ();
 sg13g2_decap_4 FILLER_86_631 ();
 sg13g2_fill_2 FILLER_86_658 ();
 sg13g2_fill_1 FILLER_86_665 ();
 sg13g2_fill_2 FILLER_86_708 ();
 sg13g2_fill_1 FILLER_86_734 ();
 sg13g2_decap_4 FILLER_86_745 ();
 sg13g2_fill_1 FILLER_86_749 ();
 sg13g2_fill_2 FILLER_86_765 ();
 sg13g2_fill_1 FILLER_86_767 ();
 sg13g2_fill_1 FILLER_86_777 ();
 sg13g2_decap_8 FILLER_86_797 ();
 sg13g2_fill_1 FILLER_86_804 ();
 sg13g2_decap_8 FILLER_86_846 ();
 sg13g2_decap_8 FILLER_86_853 ();
 sg13g2_decap_8 FILLER_86_860 ();
 sg13g2_decap_8 FILLER_86_867 ();
 sg13g2_decap_8 FILLER_86_874 ();
 sg13g2_decap_8 FILLER_86_881 ();
 sg13g2_decap_8 FILLER_86_888 ();
 sg13g2_decap_8 FILLER_86_895 ();
 sg13g2_decap_8 FILLER_86_902 ();
 sg13g2_decap_8 FILLER_86_909 ();
 sg13g2_decap_8 FILLER_86_916 ();
 sg13g2_decap_8 FILLER_86_923 ();
 sg13g2_decap_8 FILLER_86_930 ();
 sg13g2_decap_8 FILLER_86_937 ();
 sg13g2_decap_8 FILLER_86_944 ();
 sg13g2_decap_8 FILLER_86_951 ();
 sg13g2_decap_8 FILLER_86_958 ();
 sg13g2_decap_8 FILLER_86_965 ();
 sg13g2_decap_8 FILLER_86_972 ();
 sg13g2_decap_8 FILLER_86_979 ();
 sg13g2_decap_8 FILLER_86_986 ();
 sg13g2_decap_8 FILLER_86_993 ();
 sg13g2_decap_8 FILLER_86_1000 ();
 sg13g2_decap_8 FILLER_86_1007 ();
 sg13g2_decap_8 FILLER_86_1014 ();
 sg13g2_decap_8 FILLER_86_1021 ();
 sg13g2_fill_1 FILLER_86_1028 ();
 sg13g2_fill_2 FILLER_87_80 ();
 sg13g2_fill_1 FILLER_87_101 ();
 sg13g2_fill_2 FILLER_87_163 ();
 sg13g2_fill_1 FILLER_87_165 ();
 sg13g2_fill_2 FILLER_87_176 ();
 sg13g2_fill_1 FILLER_87_178 ();
 sg13g2_decap_4 FILLER_87_252 ();
 sg13g2_fill_2 FILLER_87_256 ();
 sg13g2_decap_8 FILLER_87_277 ();
 sg13g2_decap_8 FILLER_87_284 ();
 sg13g2_fill_2 FILLER_87_291 ();
 sg13g2_decap_4 FILLER_87_321 ();
 sg13g2_fill_2 FILLER_87_333 ();
 sg13g2_fill_1 FILLER_87_335 ();
 sg13g2_fill_2 FILLER_87_344 ();
 sg13g2_fill_1 FILLER_87_360 ();
 sg13g2_decap_4 FILLER_87_386 ();
 sg13g2_decap_8 FILLER_87_407 ();
 sg13g2_fill_2 FILLER_87_420 ();
 sg13g2_decap_4 FILLER_87_442 ();
 sg13g2_fill_1 FILLER_87_446 ();
 sg13g2_fill_2 FILLER_87_473 ();
 sg13g2_fill_1 FILLER_87_475 ();
 sg13g2_fill_2 FILLER_87_484 ();
 sg13g2_fill_1 FILLER_87_486 ();
 sg13g2_fill_2 FILLER_87_500 ();
 sg13g2_fill_1 FILLER_87_502 ();
 sg13g2_fill_1 FILLER_87_506 ();
 sg13g2_decap_8 FILLER_87_511 ();
 sg13g2_fill_2 FILLER_87_518 ();
 sg13g2_fill_1 FILLER_87_520 ();
 sg13g2_fill_1 FILLER_87_536 ();
 sg13g2_fill_1 FILLER_87_567 ();
 sg13g2_decap_8 FILLER_87_576 ();
 sg13g2_decap_4 FILLER_87_583 ();
 sg13g2_decap_8 FILLER_87_592 ();
 sg13g2_fill_2 FILLER_87_610 ();
 sg13g2_decap_8 FILLER_87_633 ();
 sg13g2_fill_2 FILLER_87_640 ();
 sg13g2_fill_1 FILLER_87_642 ();
 sg13g2_fill_1 FILLER_87_649 ();
 sg13g2_fill_2 FILLER_87_659 ();
 sg13g2_fill_2 FILLER_87_669 ();
 sg13g2_decap_4 FILLER_87_684 ();
 sg13g2_fill_1 FILLER_87_688 ();
 sg13g2_fill_2 FILLER_87_704 ();
 sg13g2_fill_2 FILLER_87_710 ();
 sg13g2_decap_4 FILLER_87_728 ();
 sg13g2_decap_8 FILLER_87_741 ();
 sg13g2_decap_4 FILLER_87_748 ();
 sg13g2_fill_2 FILLER_87_762 ();
 sg13g2_fill_1 FILLER_87_768 ();
 sg13g2_decap_4 FILLER_87_778 ();
 sg13g2_fill_2 FILLER_87_782 ();
 sg13g2_decap_8 FILLER_87_788 ();
 sg13g2_fill_1 FILLER_87_795 ();
 sg13g2_decap_8 FILLER_87_804 ();
 sg13g2_decap_8 FILLER_87_853 ();
 sg13g2_decap_8 FILLER_87_860 ();
 sg13g2_decap_8 FILLER_87_867 ();
 sg13g2_decap_8 FILLER_87_874 ();
 sg13g2_decap_8 FILLER_87_881 ();
 sg13g2_decap_8 FILLER_87_888 ();
 sg13g2_decap_8 FILLER_87_895 ();
 sg13g2_decap_8 FILLER_87_902 ();
 sg13g2_decap_8 FILLER_87_909 ();
 sg13g2_decap_8 FILLER_87_916 ();
 sg13g2_decap_8 FILLER_87_923 ();
 sg13g2_decap_8 FILLER_87_930 ();
 sg13g2_decap_8 FILLER_87_937 ();
 sg13g2_decap_8 FILLER_87_944 ();
 sg13g2_decap_8 FILLER_87_951 ();
 sg13g2_decap_8 FILLER_87_958 ();
 sg13g2_decap_8 FILLER_87_965 ();
 sg13g2_decap_8 FILLER_87_972 ();
 sg13g2_decap_8 FILLER_87_979 ();
 sg13g2_decap_8 FILLER_87_986 ();
 sg13g2_decap_8 FILLER_87_993 ();
 sg13g2_decap_8 FILLER_87_1000 ();
 sg13g2_decap_8 FILLER_87_1007 ();
 sg13g2_decap_8 FILLER_87_1014 ();
 sg13g2_decap_8 FILLER_87_1021 ();
 sg13g2_fill_1 FILLER_87_1028 ();
 sg13g2_fill_2 FILLER_88_0 ();
 sg13g2_decap_4 FILLER_88_17 ();
 sg13g2_decap_4 FILLER_88_30 ();
 sg13g2_decap_8 FILLER_88_43 ();
 sg13g2_decap_4 FILLER_88_143 ();
 sg13g2_fill_1 FILLER_88_147 ();
 sg13g2_decap_4 FILLER_88_175 ();
 sg13g2_fill_2 FILLER_88_179 ();
 sg13g2_decap_4 FILLER_88_200 ();
 sg13g2_fill_2 FILLER_88_227 ();
 sg13g2_fill_1 FILLER_88_229 ();
 sg13g2_decap_4 FILLER_88_249 ();
 sg13g2_fill_2 FILLER_88_253 ();
 sg13g2_fill_2 FILLER_88_281 ();
 sg13g2_fill_1 FILLER_88_301 ();
 sg13g2_fill_2 FILLER_88_316 ();
 sg13g2_fill_1 FILLER_88_318 ();
 sg13g2_fill_2 FILLER_88_343 ();
 sg13g2_fill_1 FILLER_88_345 ();
 sg13g2_fill_2 FILLER_88_354 ();
 sg13g2_decap_4 FILLER_88_362 ();
 sg13g2_fill_2 FILLER_88_387 ();
 sg13g2_decap_8 FILLER_88_400 ();
 sg13g2_decap_8 FILLER_88_407 ();
 sg13g2_fill_2 FILLER_88_414 ();
 sg13g2_fill_1 FILLER_88_416 ();
 sg13g2_decap_4 FILLER_88_430 ();
 sg13g2_fill_1 FILLER_88_434 ();
 sg13g2_fill_1 FILLER_88_440 ();
 sg13g2_decap_4 FILLER_88_446 ();
 sg13g2_fill_1 FILLER_88_450 ();
 sg13g2_fill_2 FILLER_88_456 ();
 sg13g2_fill_1 FILLER_88_458 ();
 sg13g2_decap_8 FILLER_88_465 ();
 sg13g2_decap_4 FILLER_88_472 ();
 sg13g2_fill_1 FILLER_88_476 ();
 sg13g2_fill_1 FILLER_88_503 ();
 sg13g2_decap_8 FILLER_88_509 ();
 sg13g2_decap_4 FILLER_88_516 ();
 sg13g2_fill_1 FILLER_88_529 ();
 sg13g2_decap_8 FILLER_88_540 ();
 sg13g2_fill_2 FILLER_88_562 ();
 sg13g2_decap_4 FILLER_88_571 ();
 sg13g2_fill_2 FILLER_88_575 ();
 sg13g2_decap_8 FILLER_88_585 ();
 sg13g2_decap_8 FILLER_88_592 ();
 sg13g2_decap_8 FILLER_88_603 ();
 sg13g2_decap_8 FILLER_88_610 ();
 sg13g2_decap_8 FILLER_88_617 ();
 sg13g2_decap_4 FILLER_88_624 ();
 sg13g2_decap_8 FILLER_88_641 ();
 sg13g2_decap_8 FILLER_88_648 ();
 sg13g2_decap_8 FILLER_88_658 ();
 sg13g2_decap_8 FILLER_88_665 ();
 sg13g2_decap_4 FILLER_88_689 ();
 sg13g2_fill_1 FILLER_88_693 ();
 sg13g2_decap_8 FILLER_88_699 ();
 sg13g2_decap_8 FILLER_88_706 ();
 sg13g2_decap_8 FILLER_88_713 ();
 sg13g2_decap_8 FILLER_88_720 ();
 sg13g2_fill_2 FILLER_88_727 ();
 sg13g2_fill_1 FILLER_88_729 ();
 sg13g2_fill_1 FILLER_88_734 ();
 sg13g2_decap_8 FILLER_88_751 ();
 sg13g2_fill_1 FILLER_88_778 ();
 sg13g2_fill_2 FILLER_88_788 ();
 sg13g2_decap_8 FILLER_88_808 ();
 sg13g2_decap_8 FILLER_88_815 ();
 sg13g2_decap_8 FILLER_88_847 ();
 sg13g2_decap_8 FILLER_88_854 ();
 sg13g2_decap_8 FILLER_88_861 ();
 sg13g2_decap_8 FILLER_88_868 ();
 sg13g2_decap_8 FILLER_88_875 ();
 sg13g2_decap_8 FILLER_88_882 ();
 sg13g2_decap_8 FILLER_88_889 ();
 sg13g2_decap_8 FILLER_88_896 ();
 sg13g2_decap_8 FILLER_88_903 ();
 sg13g2_decap_8 FILLER_88_910 ();
 sg13g2_decap_8 FILLER_88_917 ();
 sg13g2_decap_8 FILLER_88_924 ();
 sg13g2_decap_8 FILLER_88_931 ();
 sg13g2_decap_8 FILLER_88_938 ();
 sg13g2_decap_8 FILLER_88_945 ();
 sg13g2_decap_8 FILLER_88_952 ();
 sg13g2_decap_8 FILLER_88_959 ();
 sg13g2_decap_8 FILLER_88_966 ();
 sg13g2_decap_8 FILLER_88_973 ();
 sg13g2_decap_8 FILLER_88_980 ();
 sg13g2_decap_8 FILLER_88_987 ();
 sg13g2_decap_8 FILLER_88_994 ();
 sg13g2_decap_8 FILLER_88_1001 ();
 sg13g2_decap_8 FILLER_88_1008 ();
 sg13g2_decap_8 FILLER_88_1015 ();
 sg13g2_decap_8 FILLER_88_1022 ();
 sg13g2_fill_2 FILLER_89_93 ();
 sg13g2_decap_8 FILLER_89_153 ();
 sg13g2_fill_1 FILLER_89_160 ();
 sg13g2_decap_8 FILLER_89_207 ();
 sg13g2_fill_1 FILLER_89_214 ();
 sg13g2_decap_4 FILLER_89_332 ();
 sg13g2_fill_1 FILLER_89_336 ();
 sg13g2_decap_8 FILLER_89_348 ();
 sg13g2_decap_8 FILLER_89_355 ();
 sg13g2_fill_2 FILLER_89_362 ();
 sg13g2_fill_1 FILLER_89_364 ();
 sg13g2_decap_8 FILLER_89_371 ();
 sg13g2_fill_1 FILLER_89_378 ();
 sg13g2_fill_2 FILLER_89_383 ();
 sg13g2_decap_8 FILLER_89_398 ();
 sg13g2_decap_4 FILLER_89_405 ();
 sg13g2_fill_1 FILLER_89_409 ();
 sg13g2_fill_2 FILLER_89_438 ();
 sg13g2_fill_1 FILLER_89_440 ();
 sg13g2_fill_1 FILLER_89_451 ();
 sg13g2_fill_1 FILLER_89_459 ();
 sg13g2_fill_1 FILLER_89_473 ();
 sg13g2_fill_1 FILLER_89_482 ();
 sg13g2_fill_2 FILLER_89_496 ();
 sg13g2_fill_1 FILLER_89_498 ();
 sg13g2_fill_2 FILLER_89_519 ();
 sg13g2_decap_8 FILLER_89_539 ();
 sg13g2_decap_8 FILLER_89_546 ();
 sg13g2_decap_4 FILLER_89_553 ();
 sg13g2_fill_2 FILLER_89_557 ();
 sg13g2_decap_8 FILLER_89_565 ();
 sg13g2_decap_8 FILLER_89_572 ();
 sg13g2_fill_1 FILLER_89_579 ();
 sg13g2_fill_1 FILLER_89_585 ();
 sg13g2_fill_2 FILLER_89_595 ();
 sg13g2_fill_1 FILLER_89_610 ();
 sg13g2_decap_4 FILLER_89_618 ();
 sg13g2_fill_2 FILLER_89_622 ();
 sg13g2_fill_1 FILLER_89_635 ();
 sg13g2_decap_4 FILLER_89_640 ();
 sg13g2_fill_2 FILLER_89_644 ();
 sg13g2_fill_2 FILLER_89_656 ();
 sg13g2_decap_8 FILLER_89_664 ();
 sg13g2_decap_8 FILLER_89_671 ();
 sg13g2_decap_4 FILLER_89_678 ();
 sg13g2_fill_2 FILLER_89_682 ();
 sg13g2_fill_2 FILLER_89_689 ();
 sg13g2_fill_1 FILLER_89_691 ();
 sg13g2_decap_8 FILLER_89_706 ();
 sg13g2_fill_2 FILLER_89_713 ();
 sg13g2_fill_1 FILLER_89_715 ();
 sg13g2_fill_2 FILLER_89_727 ();
 sg13g2_fill_1 FILLER_89_729 ();
 sg13g2_fill_1 FILLER_89_742 ();
 sg13g2_decap_8 FILLER_89_758 ();
 sg13g2_decap_4 FILLER_89_765 ();
 sg13g2_fill_1 FILLER_89_790 ();
 sg13g2_decap_8 FILLER_89_811 ();
 sg13g2_decap_8 FILLER_89_818 ();
 sg13g2_decap_8 FILLER_89_839 ();
 sg13g2_decap_8 FILLER_89_846 ();
 sg13g2_decap_8 FILLER_89_853 ();
 sg13g2_decap_8 FILLER_89_860 ();
 sg13g2_decap_8 FILLER_89_867 ();
 sg13g2_decap_8 FILLER_89_874 ();
 sg13g2_decap_8 FILLER_89_881 ();
 sg13g2_decap_8 FILLER_89_888 ();
 sg13g2_decap_8 FILLER_89_895 ();
 sg13g2_decap_8 FILLER_89_902 ();
 sg13g2_decap_8 FILLER_89_909 ();
 sg13g2_decap_8 FILLER_89_916 ();
 sg13g2_decap_8 FILLER_89_923 ();
 sg13g2_decap_8 FILLER_89_930 ();
 sg13g2_decap_8 FILLER_89_937 ();
 sg13g2_decap_8 FILLER_89_944 ();
 sg13g2_decap_8 FILLER_89_951 ();
 sg13g2_decap_8 FILLER_89_958 ();
 sg13g2_decap_8 FILLER_89_965 ();
 sg13g2_decap_8 FILLER_89_972 ();
 sg13g2_decap_8 FILLER_89_979 ();
 sg13g2_decap_8 FILLER_89_986 ();
 sg13g2_decap_8 FILLER_89_993 ();
 sg13g2_decap_8 FILLER_89_1000 ();
 sg13g2_decap_8 FILLER_89_1007 ();
 sg13g2_decap_8 FILLER_89_1014 ();
 sg13g2_decap_8 FILLER_89_1021 ();
 sg13g2_fill_1 FILLER_89_1028 ();
 sg13g2_decap_8 FILLER_90_0 ();
 sg13g2_decap_8 FILLER_90_7 ();
 sg13g2_decap_8 FILLER_90_14 ();
 sg13g2_decap_8 FILLER_90_21 ();
 sg13g2_decap_8 FILLER_90_28 ();
 sg13g2_fill_1 FILLER_90_38 ();
 sg13g2_decap_4 FILLER_90_126 ();
 sg13g2_fill_2 FILLER_90_130 ();
 sg13g2_fill_2 FILLER_90_159 ();
 sg13g2_decap_4 FILLER_90_180 ();
 sg13g2_decap_4 FILLER_90_194 ();
 sg13g2_fill_2 FILLER_90_198 ();
 sg13g2_decap_4 FILLER_90_240 ();
 sg13g2_fill_1 FILLER_90_244 ();
 sg13g2_fill_2 FILLER_90_270 ();
 sg13g2_fill_1 FILLER_90_278 ();
 sg13g2_fill_2 FILLER_90_295 ();
 sg13g2_decap_8 FILLER_90_350 ();
 sg13g2_decap_8 FILLER_90_357 ();
 sg13g2_decap_4 FILLER_90_364 ();
 sg13g2_fill_1 FILLER_90_368 ();
 sg13g2_fill_2 FILLER_90_373 ();
 sg13g2_fill_1 FILLER_90_380 ();
 sg13g2_fill_2 FILLER_90_393 ();
 sg13g2_decap_8 FILLER_90_407 ();
 sg13g2_fill_1 FILLER_90_422 ();
 sg13g2_decap_8 FILLER_90_433 ();
 sg13g2_fill_1 FILLER_90_440 ();
 sg13g2_decap_8 FILLER_90_445 ();
 sg13g2_decap_8 FILLER_90_452 ();
 sg13g2_decap_8 FILLER_90_459 ();
 sg13g2_decap_8 FILLER_90_466 ();
 sg13g2_fill_2 FILLER_90_473 ();
 sg13g2_fill_1 FILLER_90_475 ();
 sg13g2_decap_8 FILLER_90_482 ();
 sg13g2_decap_8 FILLER_90_489 ();
 sg13g2_fill_2 FILLER_90_496 ();
 sg13g2_decap_8 FILLER_90_503 ();
 sg13g2_decap_8 FILLER_90_510 ();
 sg13g2_decap_4 FILLER_90_517 ();
 sg13g2_fill_2 FILLER_90_547 ();
 sg13g2_fill_1 FILLER_90_549 ();
 sg13g2_decap_4 FILLER_90_568 ();
 sg13g2_fill_2 FILLER_90_572 ();
 sg13g2_decap_4 FILLER_90_613 ();
 sg13g2_decap_8 FILLER_90_666 ();
 sg13g2_fill_2 FILLER_90_678 ();
 sg13g2_fill_1 FILLER_90_680 ();
 sg13g2_fill_2 FILLER_90_686 ();
 sg13g2_decap_8 FILLER_90_718 ();
 sg13g2_decap_8 FILLER_90_729 ();
 sg13g2_fill_2 FILLER_90_736 ();
 sg13g2_fill_1 FILLER_90_738 ();
 sg13g2_fill_2 FILLER_90_763 ();
 sg13g2_decap_4 FILLER_90_799 ();
 sg13g2_fill_2 FILLER_90_803 ();
 sg13g2_decap_8 FILLER_90_813 ();
 sg13g2_decap_8 FILLER_90_840 ();
 sg13g2_decap_8 FILLER_90_847 ();
 sg13g2_decap_8 FILLER_90_854 ();
 sg13g2_decap_8 FILLER_90_861 ();
 sg13g2_decap_8 FILLER_90_868 ();
 sg13g2_decap_8 FILLER_90_875 ();
 sg13g2_decap_8 FILLER_90_882 ();
 sg13g2_decap_8 FILLER_90_889 ();
 sg13g2_decap_8 FILLER_90_896 ();
 sg13g2_decap_8 FILLER_90_903 ();
 sg13g2_decap_8 FILLER_90_910 ();
 sg13g2_decap_8 FILLER_90_917 ();
 sg13g2_decap_8 FILLER_90_924 ();
 sg13g2_decap_8 FILLER_90_931 ();
 sg13g2_decap_8 FILLER_90_938 ();
 sg13g2_decap_8 FILLER_90_945 ();
 sg13g2_decap_8 FILLER_90_952 ();
 sg13g2_decap_8 FILLER_90_959 ();
 sg13g2_decap_8 FILLER_90_966 ();
 sg13g2_decap_8 FILLER_90_973 ();
 sg13g2_decap_8 FILLER_90_980 ();
 sg13g2_decap_8 FILLER_90_987 ();
 sg13g2_decap_8 FILLER_90_994 ();
 sg13g2_decap_8 FILLER_90_1001 ();
 sg13g2_decap_8 FILLER_90_1008 ();
 sg13g2_decap_8 FILLER_90_1015 ();
 sg13g2_decap_8 FILLER_90_1022 ();
 sg13g2_decap_8 FILLER_91_0 ();
 sg13g2_decap_8 FILLER_91_7 ();
 sg13g2_decap_8 FILLER_91_14 ();
 sg13g2_decap_8 FILLER_91_21 ();
 sg13g2_decap_4 FILLER_91_28 ();
 sg13g2_fill_1 FILLER_91_32 ();
 sg13g2_fill_2 FILLER_91_67 ();
 sg13g2_decap_4 FILLER_91_198 ();
 sg13g2_fill_2 FILLER_91_202 ();
 sg13g2_fill_2 FILLER_91_281 ();
 sg13g2_fill_2 FILLER_91_305 ();
 sg13g2_decap_8 FILLER_91_316 ();
 sg13g2_fill_2 FILLER_91_323 ();
 sg13g2_fill_1 FILLER_91_325 ();
 sg13g2_fill_1 FILLER_91_362 ();
 sg13g2_decap_8 FILLER_91_410 ();
 sg13g2_fill_1 FILLER_91_417 ();
 sg13g2_decap_8 FILLER_91_427 ();
 sg13g2_decap_8 FILLER_91_434 ();
 sg13g2_decap_4 FILLER_91_441 ();
 sg13g2_fill_1 FILLER_91_466 ();
 sg13g2_fill_1 FILLER_91_476 ();
 sg13g2_fill_2 FILLER_91_488 ();
 sg13g2_decap_8 FILLER_91_515 ();
 sg13g2_fill_2 FILLER_91_534 ();
 sg13g2_fill_2 FILLER_91_548 ();
 sg13g2_fill_1 FILLER_91_550 ();
 sg13g2_fill_2 FILLER_91_556 ();
 sg13g2_decap_8 FILLER_91_562 ();
 sg13g2_fill_1 FILLER_91_569 ();
 sg13g2_decap_4 FILLER_91_580 ();
 sg13g2_fill_2 FILLER_91_584 ();
 sg13g2_decap_4 FILLER_91_592 ();
 sg13g2_fill_1 FILLER_91_601 ();
 sg13g2_decap_4 FILLER_91_639 ();
 sg13g2_fill_2 FILLER_91_666 ();
 sg13g2_fill_2 FILLER_91_677 ();
 sg13g2_fill_1 FILLER_91_679 ();
 sg13g2_fill_1 FILLER_91_688 ();
 sg13g2_fill_1 FILLER_91_698 ();
 sg13g2_fill_1 FILLER_91_704 ();
 sg13g2_fill_2 FILLER_91_731 ();
 sg13g2_decap_8 FILLER_91_737 ();
 sg13g2_fill_2 FILLER_91_744 ();
 sg13g2_fill_1 FILLER_91_746 ();
 sg13g2_decap_8 FILLER_91_761 ();
 sg13g2_decap_8 FILLER_91_768 ();
 sg13g2_decap_8 FILLER_91_797 ();
 sg13g2_decap_4 FILLER_91_804 ();
 sg13g2_decap_8 FILLER_91_842 ();
 sg13g2_decap_8 FILLER_91_849 ();
 sg13g2_decap_8 FILLER_91_856 ();
 sg13g2_decap_8 FILLER_91_863 ();
 sg13g2_decap_8 FILLER_91_870 ();
 sg13g2_decap_8 FILLER_91_877 ();
 sg13g2_decap_8 FILLER_91_884 ();
 sg13g2_decap_8 FILLER_91_891 ();
 sg13g2_decap_8 FILLER_91_898 ();
 sg13g2_decap_8 FILLER_91_905 ();
 sg13g2_decap_8 FILLER_91_912 ();
 sg13g2_decap_8 FILLER_91_919 ();
 sg13g2_decap_8 FILLER_91_926 ();
 sg13g2_decap_8 FILLER_91_933 ();
 sg13g2_decap_8 FILLER_91_940 ();
 sg13g2_decap_8 FILLER_91_947 ();
 sg13g2_decap_8 FILLER_91_954 ();
 sg13g2_decap_8 FILLER_91_961 ();
 sg13g2_decap_8 FILLER_91_968 ();
 sg13g2_decap_8 FILLER_91_975 ();
 sg13g2_decap_8 FILLER_91_982 ();
 sg13g2_decap_8 FILLER_91_989 ();
 sg13g2_decap_8 FILLER_91_996 ();
 sg13g2_decap_8 FILLER_91_1003 ();
 sg13g2_decap_8 FILLER_91_1010 ();
 sg13g2_decap_8 FILLER_91_1017 ();
 sg13g2_decap_4 FILLER_91_1024 ();
 sg13g2_fill_1 FILLER_91_1028 ();
 sg13g2_decap_8 FILLER_92_0 ();
 sg13g2_decap_8 FILLER_92_7 ();
 sg13g2_decap_8 FILLER_92_14 ();
 sg13g2_decap_8 FILLER_92_21 ();
 sg13g2_decap_8 FILLER_92_28 ();
 sg13g2_decap_4 FILLER_92_35 ();
 sg13g2_fill_1 FILLER_92_67 ();
 sg13g2_fill_2 FILLER_92_132 ();
 sg13g2_decap_8 FILLER_92_144 ();
 sg13g2_decap_8 FILLER_92_160 ();
 sg13g2_fill_1 FILLER_92_167 ();
 sg13g2_fill_2 FILLER_92_278 ();
 sg13g2_fill_1 FILLER_92_293 ();
 sg13g2_decap_8 FILLER_92_319 ();
 sg13g2_decap_4 FILLER_92_326 ();
 sg13g2_fill_1 FILLER_92_335 ();
 sg13g2_decap_4 FILLER_92_341 ();
 sg13g2_fill_2 FILLER_92_345 ();
 sg13g2_fill_2 FILLER_92_352 ();
 sg13g2_decap_4 FILLER_92_362 ();
 sg13g2_fill_1 FILLER_92_366 ();
 sg13g2_fill_1 FILLER_92_373 ();
 sg13g2_fill_2 FILLER_92_382 ();
 sg13g2_decap_8 FILLER_92_400 ();
 sg13g2_decap_4 FILLER_92_407 ();
 sg13g2_fill_2 FILLER_92_436 ();
 sg13g2_fill_1 FILLER_92_438 ();
 sg13g2_fill_1 FILLER_92_449 ();
 sg13g2_decap_8 FILLER_92_464 ();
 sg13g2_decap_8 FILLER_92_471 ();
 sg13g2_fill_1 FILLER_92_503 ();
 sg13g2_decap_8 FILLER_92_527 ();
 sg13g2_decap_4 FILLER_92_534 ();
 sg13g2_fill_2 FILLER_92_538 ();
 sg13g2_fill_2 FILLER_92_545 ();
 sg13g2_fill_1 FILLER_92_552 ();
 sg13g2_fill_2 FILLER_92_569 ();
 sg13g2_fill_1 FILLER_92_571 ();
 sg13g2_fill_1 FILLER_92_585 ();
 sg13g2_fill_2 FILLER_92_599 ();
 sg13g2_fill_1 FILLER_92_601 ();
 sg13g2_decap_8 FILLER_92_606 ();
 sg13g2_fill_2 FILLER_92_613 ();
 sg13g2_fill_2 FILLER_92_619 ();
 sg13g2_decap_4 FILLER_92_641 ();
 sg13g2_decap_8 FILLER_92_648 ();
 sg13g2_fill_1 FILLER_92_664 ();
 sg13g2_decap_8 FILLER_92_670 ();
 sg13g2_fill_2 FILLER_92_677 ();
 sg13g2_fill_1 FILLER_92_679 ();
 sg13g2_decap_4 FILLER_92_684 ();
 sg13g2_fill_2 FILLER_92_696 ();
 sg13g2_fill_1 FILLER_92_698 ();
 sg13g2_decap_4 FILLER_92_704 ();
 sg13g2_fill_2 FILLER_92_708 ();
 sg13g2_fill_2 FILLER_92_721 ();
 sg13g2_fill_2 FILLER_92_738 ();
 sg13g2_fill_1 FILLER_92_740 ();
 sg13g2_decap_4 FILLER_92_746 ();
 sg13g2_fill_1 FILLER_92_750 ();
 sg13g2_decap_8 FILLER_92_755 ();
 sg13g2_decap_8 FILLER_92_762 ();
 sg13g2_fill_2 FILLER_92_769 ();
 sg13g2_fill_1 FILLER_92_771 ();
 sg13g2_decap_8 FILLER_92_789 ();
 sg13g2_fill_2 FILLER_92_796 ();
 sg13g2_decap_8 FILLER_92_806 ();
 sg13g2_decap_4 FILLER_92_813 ();
 sg13g2_fill_2 FILLER_92_817 ();
 sg13g2_decap_8 FILLER_92_836 ();
 sg13g2_decap_8 FILLER_92_843 ();
 sg13g2_decap_8 FILLER_92_850 ();
 sg13g2_decap_8 FILLER_92_857 ();
 sg13g2_decap_8 FILLER_92_864 ();
 sg13g2_decap_8 FILLER_92_871 ();
 sg13g2_decap_8 FILLER_92_878 ();
 sg13g2_decap_8 FILLER_92_885 ();
 sg13g2_decap_8 FILLER_92_892 ();
 sg13g2_decap_8 FILLER_92_899 ();
 sg13g2_decap_8 FILLER_92_906 ();
 sg13g2_decap_8 FILLER_92_913 ();
 sg13g2_decap_8 FILLER_92_920 ();
 sg13g2_decap_8 FILLER_92_927 ();
 sg13g2_decap_8 FILLER_92_934 ();
 sg13g2_decap_8 FILLER_92_941 ();
 sg13g2_decap_8 FILLER_92_948 ();
 sg13g2_decap_8 FILLER_92_955 ();
 sg13g2_decap_8 FILLER_92_962 ();
 sg13g2_decap_8 FILLER_92_969 ();
 sg13g2_decap_8 FILLER_92_976 ();
 sg13g2_decap_8 FILLER_92_983 ();
 sg13g2_decap_8 FILLER_92_990 ();
 sg13g2_decap_8 FILLER_92_997 ();
 sg13g2_decap_8 FILLER_92_1004 ();
 sg13g2_decap_8 FILLER_92_1011 ();
 sg13g2_decap_8 FILLER_92_1018 ();
 sg13g2_decap_4 FILLER_92_1025 ();
 sg13g2_decap_8 FILLER_93_0 ();
 sg13g2_decap_8 FILLER_93_7 ();
 sg13g2_decap_8 FILLER_93_14 ();
 sg13g2_decap_8 FILLER_93_21 ();
 sg13g2_decap_8 FILLER_93_28 ();
 sg13g2_decap_8 FILLER_93_35 ();
 sg13g2_decap_8 FILLER_93_42 ();
 sg13g2_fill_2 FILLER_93_49 ();
 sg13g2_fill_1 FILLER_93_51 ();
 sg13g2_decap_8 FILLER_93_92 ();
 sg13g2_decap_8 FILLER_93_112 ();
 sg13g2_fill_1 FILLER_93_129 ();
 sg13g2_fill_2 FILLER_93_177 ();
 sg13g2_fill_1 FILLER_93_179 ();
 sg13g2_decap_4 FILLER_93_190 ();
 sg13g2_fill_2 FILLER_93_194 ();
 sg13g2_decap_4 FILLER_93_209 ();
 sg13g2_fill_2 FILLER_93_213 ();
 sg13g2_fill_2 FILLER_93_250 ();
 sg13g2_fill_1 FILLER_93_252 ();
 sg13g2_fill_1 FILLER_93_262 ();
 sg13g2_decap_4 FILLER_93_293 ();
 sg13g2_fill_1 FILLER_93_297 ();
 sg13g2_fill_1 FILLER_93_303 ();
 sg13g2_fill_2 FILLER_93_319 ();
 sg13g2_fill_1 FILLER_93_321 ();
 sg13g2_fill_1 FILLER_93_330 ();
 sg13g2_fill_2 FILLER_93_352 ();
 sg13g2_fill_1 FILLER_93_354 ();
 sg13g2_fill_2 FILLER_93_366 ();
 sg13g2_fill_1 FILLER_93_368 ();
 sg13g2_decap_8 FILLER_93_400 ();
 sg13g2_decap_8 FILLER_93_407 ();
 sg13g2_decap_8 FILLER_93_414 ();
 sg13g2_fill_2 FILLER_93_434 ();
 sg13g2_fill_1 FILLER_93_436 ();
 sg13g2_fill_2 FILLER_93_452 ();
 sg13g2_decap_4 FILLER_93_459 ();
 sg13g2_fill_1 FILLER_93_463 ();
 sg13g2_decap_8 FILLER_93_495 ();
 sg13g2_decap_8 FILLER_93_502 ();
 sg13g2_decap_8 FILLER_93_509 ();
 sg13g2_decap_8 FILLER_93_516 ();
 sg13g2_fill_2 FILLER_93_523 ();
 sg13g2_decap_8 FILLER_93_537 ();
 sg13g2_fill_2 FILLER_93_544 ();
 sg13g2_fill_1 FILLER_93_554 ();
 sg13g2_decap_8 FILLER_93_560 ();
 sg13g2_decap_4 FILLER_93_567 ();
 sg13g2_fill_1 FILLER_93_571 ();
 sg13g2_fill_2 FILLER_93_624 ();
 sg13g2_fill_2 FILLER_93_639 ();
 sg13g2_decap_4 FILLER_93_649 ();
 sg13g2_fill_2 FILLER_93_653 ();
 sg13g2_decap_8 FILLER_93_673 ();
 sg13g2_fill_2 FILLER_93_708 ();
 sg13g2_fill_1 FILLER_93_710 ();
 sg13g2_fill_2 FILLER_93_716 ();
 sg13g2_fill_1 FILLER_93_718 ();
 sg13g2_decap_8 FILLER_93_729 ();
 sg13g2_fill_2 FILLER_93_736 ();
 sg13g2_decap_4 FILLER_93_742 ();
 sg13g2_fill_2 FILLER_93_746 ();
 sg13g2_decap_8 FILLER_93_754 ();
 sg13g2_fill_1 FILLER_93_761 ();
 sg13g2_decap_8 FILLER_93_800 ();
 sg13g2_fill_1 FILLER_93_807 ();
 sg13g2_fill_1 FILLER_93_822 ();
 sg13g2_decap_8 FILLER_93_832 ();
 sg13g2_decap_8 FILLER_93_839 ();
 sg13g2_decap_8 FILLER_93_846 ();
 sg13g2_decap_8 FILLER_93_853 ();
 sg13g2_decap_8 FILLER_93_860 ();
 sg13g2_decap_8 FILLER_93_867 ();
 sg13g2_decap_8 FILLER_93_874 ();
 sg13g2_decap_8 FILLER_93_881 ();
 sg13g2_decap_8 FILLER_93_888 ();
 sg13g2_decap_8 FILLER_93_895 ();
 sg13g2_decap_8 FILLER_93_902 ();
 sg13g2_decap_8 FILLER_93_909 ();
 sg13g2_decap_8 FILLER_93_916 ();
 sg13g2_decap_8 FILLER_93_923 ();
 sg13g2_decap_8 FILLER_93_930 ();
 sg13g2_decap_8 FILLER_93_937 ();
 sg13g2_decap_8 FILLER_93_944 ();
 sg13g2_decap_8 FILLER_93_951 ();
 sg13g2_decap_8 FILLER_93_958 ();
 sg13g2_decap_8 FILLER_93_965 ();
 sg13g2_decap_8 FILLER_93_972 ();
 sg13g2_decap_8 FILLER_93_979 ();
 sg13g2_decap_8 FILLER_93_986 ();
 sg13g2_decap_8 FILLER_93_993 ();
 sg13g2_decap_8 FILLER_93_1000 ();
 sg13g2_decap_8 FILLER_93_1007 ();
 sg13g2_decap_8 FILLER_93_1014 ();
 sg13g2_decap_8 FILLER_93_1021 ();
 sg13g2_fill_1 FILLER_93_1028 ();
 sg13g2_decap_8 FILLER_94_0 ();
 sg13g2_decap_8 FILLER_94_7 ();
 sg13g2_decap_8 FILLER_94_14 ();
 sg13g2_decap_8 FILLER_94_21 ();
 sg13g2_decap_8 FILLER_94_28 ();
 sg13g2_decap_8 FILLER_94_35 ();
 sg13g2_decap_8 FILLER_94_42 ();
 sg13g2_decap_8 FILLER_94_49 ();
 sg13g2_decap_4 FILLER_94_56 ();
 sg13g2_fill_2 FILLER_94_60 ();
 sg13g2_decap_8 FILLER_94_89 ();
 sg13g2_fill_1 FILLER_94_96 ();
 sg13g2_decap_4 FILLER_94_163 ();
 sg13g2_fill_1 FILLER_94_167 ();
 sg13g2_fill_2 FILLER_94_181 ();
 sg13g2_fill_2 FILLER_94_217 ();
 sg13g2_fill_1 FILLER_94_219 ();
 sg13g2_fill_2 FILLER_94_252 ();
 sg13g2_fill_2 FILLER_94_283 ();
 sg13g2_decap_4 FILLER_94_295 ();
 sg13g2_fill_1 FILLER_94_299 ();
 sg13g2_fill_2 FILLER_94_319 ();
 sg13g2_fill_1 FILLER_94_321 ();
 sg13g2_fill_1 FILLER_94_328 ();
 sg13g2_fill_2 FILLER_94_349 ();
 sg13g2_fill_1 FILLER_94_351 ();
 sg13g2_decap_8 FILLER_94_396 ();
 sg13g2_fill_2 FILLER_94_403 ();
 sg13g2_decap_8 FILLER_94_457 ();
 sg13g2_decap_4 FILLER_94_464 ();
 sg13g2_fill_1 FILLER_94_468 ();
 sg13g2_decap_8 FILLER_94_493 ();
 sg13g2_fill_1 FILLER_94_500 ();
 sg13g2_fill_1 FILLER_94_527 ();
 sg13g2_fill_1 FILLER_94_533 ();
 sg13g2_decap_8 FILLER_94_542 ();
 sg13g2_fill_2 FILLER_94_549 ();
 sg13g2_fill_1 FILLER_94_551 ();
 sg13g2_decap_8 FILLER_94_560 ();
 sg13g2_decap_4 FILLER_94_580 ();
 sg13g2_fill_2 FILLER_94_584 ();
 sg13g2_decap_4 FILLER_94_591 ();
 sg13g2_fill_2 FILLER_94_595 ();
 sg13g2_fill_1 FILLER_94_610 ();
 sg13g2_decap_8 FILLER_94_616 ();
 sg13g2_fill_1 FILLER_94_633 ();
 sg13g2_decap_8 FILLER_94_645 ();
 sg13g2_decap_4 FILLER_94_652 ();
 sg13g2_fill_2 FILLER_94_656 ();
 sg13g2_decap_4 FILLER_94_674 ();
 sg13g2_decap_8 FILLER_94_701 ();
 sg13g2_fill_1 FILLER_94_708 ();
 sg13g2_decap_4 FILLER_94_718 ();
 sg13g2_fill_1 FILLER_94_722 ();
 sg13g2_decap_4 FILLER_94_727 ();
 sg13g2_fill_2 FILLER_94_741 ();
 sg13g2_fill_2 FILLER_94_753 ();
 sg13g2_fill_1 FILLER_94_755 ();
 sg13g2_decap_4 FILLER_94_794 ();
 sg13g2_fill_1 FILLER_94_798 ();
 sg13g2_decap_8 FILLER_94_840 ();
 sg13g2_decap_8 FILLER_94_847 ();
 sg13g2_decap_8 FILLER_94_854 ();
 sg13g2_decap_8 FILLER_94_861 ();
 sg13g2_decap_8 FILLER_94_868 ();
 sg13g2_decap_8 FILLER_94_875 ();
 sg13g2_decap_8 FILLER_94_882 ();
 sg13g2_decap_8 FILLER_94_889 ();
 sg13g2_decap_8 FILLER_94_896 ();
 sg13g2_decap_8 FILLER_94_903 ();
 sg13g2_decap_8 FILLER_94_910 ();
 sg13g2_decap_8 FILLER_94_917 ();
 sg13g2_decap_8 FILLER_94_924 ();
 sg13g2_decap_8 FILLER_94_931 ();
 sg13g2_decap_8 FILLER_94_938 ();
 sg13g2_decap_8 FILLER_94_945 ();
 sg13g2_decap_8 FILLER_94_952 ();
 sg13g2_decap_8 FILLER_94_959 ();
 sg13g2_decap_8 FILLER_94_966 ();
 sg13g2_decap_8 FILLER_94_973 ();
 sg13g2_decap_8 FILLER_94_980 ();
 sg13g2_decap_8 FILLER_94_987 ();
 sg13g2_decap_8 FILLER_94_994 ();
 sg13g2_decap_8 FILLER_94_1001 ();
 sg13g2_decap_8 FILLER_94_1008 ();
 sg13g2_decap_8 FILLER_94_1015 ();
 sg13g2_decap_8 FILLER_94_1022 ();
 sg13g2_decap_8 FILLER_95_0 ();
 sg13g2_decap_8 FILLER_95_7 ();
 sg13g2_decap_8 FILLER_95_14 ();
 sg13g2_decap_8 FILLER_95_21 ();
 sg13g2_decap_8 FILLER_95_28 ();
 sg13g2_decap_8 FILLER_95_35 ();
 sg13g2_decap_8 FILLER_95_42 ();
 sg13g2_decap_8 FILLER_95_49 ();
 sg13g2_decap_8 FILLER_95_56 ();
 sg13g2_decap_4 FILLER_95_63 ();
 sg13g2_fill_1 FILLER_95_125 ();
 sg13g2_decap_4 FILLER_95_191 ();
 sg13g2_fill_2 FILLER_95_195 ();
 sg13g2_decap_4 FILLER_95_215 ();
 sg13g2_decap_8 FILLER_95_242 ();
 sg13g2_fill_2 FILLER_95_278 ();
 sg13g2_fill_1 FILLER_95_280 ();
 sg13g2_decap_8 FILLER_95_285 ();
 sg13g2_fill_2 FILLER_95_292 ();
 sg13g2_fill_1 FILLER_95_294 ();
 sg13g2_fill_2 FILLER_95_300 ();
 sg13g2_fill_1 FILLER_95_302 ();
 sg13g2_decap_4 FILLER_95_316 ();
 sg13g2_fill_1 FILLER_95_320 ();
 sg13g2_decap_4 FILLER_95_326 ();
 sg13g2_fill_1 FILLER_95_330 ();
 sg13g2_fill_2 FILLER_95_369 ();
 sg13g2_decap_8 FILLER_95_395 ();
 sg13g2_decap_8 FILLER_95_402 ();
 sg13g2_fill_1 FILLER_95_422 ();
 sg13g2_fill_1 FILLER_95_436 ();
 sg13g2_decap_4 FILLER_95_461 ();
 sg13g2_fill_1 FILLER_95_465 ();
 sg13g2_decap_4 FILLER_95_480 ();
 sg13g2_decap_8 FILLER_95_488 ();
 sg13g2_fill_2 FILLER_95_495 ();
 sg13g2_fill_1 FILLER_95_525 ();
 sg13g2_decap_8 FILLER_95_551 ();
 sg13g2_decap_4 FILLER_95_558 ();
 sg13g2_fill_1 FILLER_95_577 ();
 sg13g2_decap_4 FILLER_95_583 ();
 sg13g2_decap_4 FILLER_95_592 ();
 sg13g2_fill_2 FILLER_95_596 ();
 sg13g2_fill_1 FILLER_95_603 ();
 sg13g2_decap_8 FILLER_95_625 ();
 sg13g2_decap_8 FILLER_95_650 ();
 sg13g2_decap_8 FILLER_95_657 ();
 sg13g2_fill_2 FILLER_95_664 ();
 sg13g2_decap_4 FILLER_95_700 ();
 sg13g2_fill_2 FILLER_95_710 ();
 sg13g2_fill_1 FILLER_95_717 ();
 sg13g2_fill_2 FILLER_95_730 ();
 sg13g2_decap_4 FILLER_95_736 ();
 sg13g2_fill_1 FILLER_95_740 ();
 sg13g2_decap_8 FILLER_95_745 ();
 sg13g2_decap_8 FILLER_95_752 ();
 sg13g2_fill_2 FILLER_95_759 ();
 sg13g2_fill_1 FILLER_95_761 ();
 sg13g2_fill_1 FILLER_95_771 ();
 sg13g2_decap_8 FILLER_95_786 ();
 sg13g2_decap_8 FILLER_95_793 ();
 sg13g2_decap_4 FILLER_95_800 ();
 sg13g2_fill_2 FILLER_95_812 ();
 sg13g2_fill_1 FILLER_95_814 ();
 sg13g2_decap_8 FILLER_95_833 ();
 sg13g2_decap_8 FILLER_95_840 ();
 sg13g2_decap_8 FILLER_95_847 ();
 sg13g2_decap_8 FILLER_95_854 ();
 sg13g2_decap_8 FILLER_95_861 ();
 sg13g2_decap_8 FILLER_95_868 ();
 sg13g2_decap_8 FILLER_95_875 ();
 sg13g2_decap_8 FILLER_95_882 ();
 sg13g2_decap_8 FILLER_95_889 ();
 sg13g2_decap_8 FILLER_95_896 ();
 sg13g2_decap_8 FILLER_95_903 ();
 sg13g2_decap_8 FILLER_95_910 ();
 sg13g2_decap_8 FILLER_95_917 ();
 sg13g2_decap_8 FILLER_95_924 ();
 sg13g2_decap_8 FILLER_95_931 ();
 sg13g2_decap_8 FILLER_95_938 ();
 sg13g2_decap_8 FILLER_95_945 ();
 sg13g2_decap_8 FILLER_95_952 ();
 sg13g2_decap_8 FILLER_95_959 ();
 sg13g2_decap_8 FILLER_95_966 ();
 sg13g2_decap_8 FILLER_95_973 ();
 sg13g2_decap_8 FILLER_95_980 ();
 sg13g2_decap_8 FILLER_95_987 ();
 sg13g2_decap_8 FILLER_95_994 ();
 sg13g2_decap_8 FILLER_95_1001 ();
 sg13g2_decap_8 FILLER_95_1008 ();
 sg13g2_decap_8 FILLER_95_1015 ();
 sg13g2_decap_8 FILLER_95_1022 ();
 sg13g2_decap_8 FILLER_96_0 ();
 sg13g2_decap_8 FILLER_96_7 ();
 sg13g2_decap_8 FILLER_96_14 ();
 sg13g2_decap_8 FILLER_96_21 ();
 sg13g2_decap_8 FILLER_96_28 ();
 sg13g2_decap_8 FILLER_96_35 ();
 sg13g2_decap_8 FILLER_96_42 ();
 sg13g2_decap_8 FILLER_96_49 ();
 sg13g2_decap_8 FILLER_96_56 ();
 sg13g2_decap_8 FILLER_96_63 ();
 sg13g2_decap_8 FILLER_96_70 ();
 sg13g2_decap_8 FILLER_96_77 ();
 sg13g2_decap_8 FILLER_96_84 ();
 sg13g2_decap_4 FILLER_96_91 ();
 sg13g2_decap_4 FILLER_96_155 ();
 sg13g2_fill_1 FILLER_96_222 ();
 sg13g2_fill_2 FILLER_96_233 ();
 sg13g2_fill_2 FILLER_96_270 ();
 sg13g2_fill_2 FILLER_96_276 ();
 sg13g2_fill_1 FILLER_96_291 ();
 sg13g2_decap_8 FILLER_96_307 ();
 sg13g2_decap_8 FILLER_96_314 ();
 sg13g2_decap_8 FILLER_96_321 ();
 sg13g2_decap_4 FILLER_96_328 ();
 sg13g2_fill_2 FILLER_96_332 ();
 sg13g2_fill_2 FILLER_96_354 ();
 sg13g2_fill_2 FILLER_96_382 ();
 sg13g2_decap_4 FILLER_96_396 ();
 sg13g2_fill_2 FILLER_96_400 ();
 sg13g2_decap_4 FILLER_96_422 ();
 sg13g2_fill_2 FILLER_96_426 ();
 sg13g2_fill_2 FILLER_96_451 ();
 sg13g2_fill_2 FILLER_96_473 ();
 sg13g2_fill_1 FILLER_96_475 ();
 sg13g2_decap_4 FILLER_96_491 ();
 sg13g2_fill_2 FILLER_96_500 ();
 sg13g2_decap_8 FILLER_96_512 ();
 sg13g2_decap_4 FILLER_96_519 ();
 sg13g2_fill_2 FILLER_96_523 ();
 sg13g2_fill_1 FILLER_96_533 ();
 sg13g2_fill_2 FILLER_96_547 ();
 sg13g2_fill_2 FILLER_96_580 ();
 sg13g2_fill_1 FILLER_96_582 ();
 sg13g2_fill_2 FILLER_96_614 ();
 sg13g2_decap_8 FILLER_96_656 ();
 sg13g2_decap_8 FILLER_96_663 ();
 sg13g2_decap_4 FILLER_96_695 ();
 sg13g2_fill_2 FILLER_96_699 ();
 sg13g2_fill_2 FILLER_96_705 ();
 sg13g2_decap_4 FILLER_96_710 ();
 sg13g2_fill_1 FILLER_96_714 ();
 sg13g2_decap_4 FILLER_96_720 ();
 sg13g2_fill_1 FILLER_96_734 ();
 sg13g2_decap_8 FILLER_96_743 ();
 sg13g2_decap_8 FILLER_96_750 ();
 sg13g2_decap_8 FILLER_96_757 ();
 sg13g2_decap_8 FILLER_96_764 ();
 sg13g2_fill_1 FILLER_96_771 ();
 sg13g2_fill_2 FILLER_96_776 ();
 sg13g2_fill_1 FILLER_96_778 ();
 sg13g2_decap_8 FILLER_96_788 ();
 sg13g2_decap_8 FILLER_96_795 ();
 sg13g2_decap_8 FILLER_96_802 ();
 sg13g2_decap_8 FILLER_96_831 ();
 sg13g2_decap_8 FILLER_96_838 ();
 sg13g2_decap_8 FILLER_96_845 ();
 sg13g2_decap_8 FILLER_96_852 ();
 sg13g2_decap_8 FILLER_96_859 ();
 sg13g2_decap_8 FILLER_96_866 ();
 sg13g2_decap_8 FILLER_96_873 ();
 sg13g2_decap_8 FILLER_96_880 ();
 sg13g2_decap_8 FILLER_96_887 ();
 sg13g2_decap_8 FILLER_96_894 ();
 sg13g2_decap_8 FILLER_96_901 ();
 sg13g2_decap_8 FILLER_96_908 ();
 sg13g2_decap_8 FILLER_96_915 ();
 sg13g2_decap_8 FILLER_96_922 ();
 sg13g2_decap_8 FILLER_96_929 ();
 sg13g2_decap_8 FILLER_96_936 ();
 sg13g2_decap_8 FILLER_96_943 ();
 sg13g2_decap_8 FILLER_96_950 ();
 sg13g2_decap_8 FILLER_96_957 ();
 sg13g2_decap_8 FILLER_96_964 ();
 sg13g2_decap_8 FILLER_96_971 ();
 sg13g2_decap_8 FILLER_96_978 ();
 sg13g2_decap_8 FILLER_96_985 ();
 sg13g2_decap_8 FILLER_96_992 ();
 sg13g2_decap_8 FILLER_96_999 ();
 sg13g2_decap_8 FILLER_96_1006 ();
 sg13g2_decap_8 FILLER_96_1013 ();
 sg13g2_decap_8 FILLER_96_1020 ();
 sg13g2_fill_2 FILLER_96_1027 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_8 FILLER_97_7 ();
 sg13g2_decap_8 FILLER_97_14 ();
 sg13g2_decap_8 FILLER_97_21 ();
 sg13g2_decap_8 FILLER_97_28 ();
 sg13g2_decap_8 FILLER_97_35 ();
 sg13g2_decap_8 FILLER_97_42 ();
 sg13g2_decap_8 FILLER_97_49 ();
 sg13g2_decap_8 FILLER_97_56 ();
 sg13g2_decap_8 FILLER_97_63 ();
 sg13g2_decap_8 FILLER_97_70 ();
 sg13g2_decap_8 FILLER_97_77 ();
 sg13g2_decap_8 FILLER_97_84 ();
 sg13g2_decap_8 FILLER_97_91 ();
 sg13g2_decap_4 FILLER_97_98 ();
 sg13g2_decap_4 FILLER_97_134 ();
 sg13g2_fill_1 FILLER_97_176 ();
 sg13g2_decap_8 FILLER_97_187 ();
 sg13g2_decap_4 FILLER_97_207 ();
 sg13g2_decap_8 FILLER_97_256 ();
 sg13g2_fill_1 FILLER_97_263 ();
 sg13g2_fill_1 FILLER_97_301 ();
 sg13g2_decap_4 FILLER_97_344 ();
 sg13g2_decap_4 FILLER_97_359 ();
 sg13g2_fill_1 FILLER_97_363 ();
 sg13g2_fill_1 FILLER_97_377 ();
 sg13g2_fill_1 FILLER_97_382 ();
 sg13g2_decap_8 FILLER_97_388 ();
 sg13g2_fill_1 FILLER_97_395 ();
 sg13g2_decap_4 FILLER_97_429 ();
 sg13g2_fill_1 FILLER_97_433 ();
 sg13g2_fill_1 FILLER_97_439 ();
 sg13g2_fill_2 FILLER_97_464 ();
 sg13g2_fill_1 FILLER_97_466 ();
 sg13g2_decap_8 FILLER_97_482 ();
 sg13g2_fill_2 FILLER_97_489 ();
 sg13g2_fill_1 FILLER_97_491 ();
 sg13g2_fill_2 FILLER_97_496 ();
 sg13g2_fill_1 FILLER_97_498 ();
 sg13g2_decap_8 FILLER_97_511 ();
 sg13g2_decap_4 FILLER_97_518 ();
 sg13g2_decap_8 FILLER_97_527 ();
 sg13g2_decap_8 FILLER_97_534 ();
 sg13g2_fill_2 FILLER_97_541 ();
 sg13g2_fill_1 FILLER_97_543 ();
 sg13g2_fill_2 FILLER_97_549 ();
 sg13g2_decap_8 FILLER_97_557 ();
 sg13g2_fill_2 FILLER_97_564 ();
 sg13g2_decap_8 FILLER_97_579 ();
 sg13g2_decap_8 FILLER_97_586 ();
 sg13g2_decap_8 FILLER_97_593 ();
 sg13g2_fill_2 FILLER_97_600 ();
 sg13g2_fill_1 FILLER_97_602 ();
 sg13g2_fill_2 FILLER_97_612 ();
 sg13g2_decap_8 FILLER_97_617 ();
 sg13g2_decap_8 FILLER_97_624 ();
 sg13g2_decap_8 FILLER_97_631 ();
 sg13g2_fill_2 FILLER_97_651 ();
 sg13g2_fill_1 FILLER_97_653 ();
 sg13g2_decap_8 FILLER_97_659 ();
 sg13g2_decap_8 FILLER_97_666 ();
 sg13g2_decap_8 FILLER_97_673 ();
 sg13g2_decap_8 FILLER_97_680 ();
 sg13g2_fill_2 FILLER_97_687 ();
 sg13g2_fill_1 FILLER_97_689 ();
 sg13g2_fill_1 FILLER_97_716 ();
 sg13g2_decap_8 FILLER_97_749 ();
 sg13g2_fill_2 FILLER_97_756 ();
 sg13g2_fill_1 FILLER_97_758 ();
 sg13g2_fill_1 FILLER_97_772 ();
 sg13g2_fill_1 FILLER_97_777 ();
 sg13g2_fill_2 FILLER_97_783 ();
 sg13g2_decap_8 FILLER_97_798 ();
 sg13g2_decap_8 FILLER_97_805 ();
 sg13g2_fill_1 FILLER_97_812 ();
 sg13g2_decap_8 FILLER_97_817 ();
 sg13g2_decap_8 FILLER_97_824 ();
 sg13g2_decap_8 FILLER_97_831 ();
 sg13g2_decap_8 FILLER_97_838 ();
 sg13g2_decap_8 FILLER_97_845 ();
 sg13g2_decap_8 FILLER_97_852 ();
 sg13g2_decap_8 FILLER_97_859 ();
 sg13g2_decap_8 FILLER_97_866 ();
 sg13g2_decap_8 FILLER_97_873 ();
 sg13g2_decap_8 FILLER_97_880 ();
 sg13g2_decap_8 FILLER_97_887 ();
 sg13g2_decap_8 FILLER_97_894 ();
 sg13g2_decap_8 FILLER_97_901 ();
 sg13g2_decap_8 FILLER_97_908 ();
 sg13g2_decap_8 FILLER_97_915 ();
 sg13g2_decap_8 FILLER_97_922 ();
 sg13g2_decap_8 FILLER_97_929 ();
 sg13g2_decap_8 FILLER_97_936 ();
 sg13g2_decap_8 FILLER_97_943 ();
 sg13g2_decap_8 FILLER_97_950 ();
 sg13g2_decap_8 FILLER_97_957 ();
 sg13g2_decap_8 FILLER_97_964 ();
 sg13g2_decap_8 FILLER_97_971 ();
 sg13g2_decap_8 FILLER_97_978 ();
 sg13g2_decap_8 FILLER_97_985 ();
 sg13g2_decap_8 FILLER_97_992 ();
 sg13g2_decap_8 FILLER_97_999 ();
 sg13g2_decap_8 FILLER_97_1006 ();
 sg13g2_decap_8 FILLER_97_1013 ();
 sg13g2_decap_8 FILLER_97_1020 ();
 sg13g2_fill_2 FILLER_97_1027 ();
 sg13g2_decap_8 FILLER_98_0 ();
 sg13g2_decap_8 FILLER_98_7 ();
 sg13g2_decap_8 FILLER_98_14 ();
 sg13g2_decap_8 FILLER_98_21 ();
 sg13g2_decap_8 FILLER_98_28 ();
 sg13g2_decap_8 FILLER_98_35 ();
 sg13g2_decap_8 FILLER_98_42 ();
 sg13g2_decap_8 FILLER_98_49 ();
 sg13g2_decap_8 FILLER_98_56 ();
 sg13g2_decap_8 FILLER_98_63 ();
 sg13g2_decap_8 FILLER_98_70 ();
 sg13g2_decap_8 FILLER_98_77 ();
 sg13g2_decap_8 FILLER_98_84 ();
 sg13g2_decap_8 FILLER_98_91 ();
 sg13g2_decap_8 FILLER_98_98 ();
 sg13g2_decap_4 FILLER_98_105 ();
 sg13g2_fill_1 FILLER_98_182 ();
 sg13g2_fill_1 FILLER_98_211 ();
 sg13g2_decap_4 FILLER_98_240 ();
 sg13g2_fill_2 FILLER_98_244 ();
 sg13g2_decap_8 FILLER_98_273 ();
 sg13g2_fill_2 FILLER_98_280 ();
 sg13g2_decap_8 FILLER_98_359 ();
 sg13g2_decap_8 FILLER_98_366 ();
 sg13g2_decap_8 FILLER_98_373 ();
 sg13g2_decap_4 FILLER_98_380 ();
 sg13g2_fill_2 FILLER_98_384 ();
 sg13g2_decap_8 FILLER_98_391 ();
 sg13g2_fill_2 FILLER_98_398 ();
 sg13g2_decap_8 FILLER_98_422 ();
 sg13g2_decap_8 FILLER_98_429 ();
 sg13g2_fill_2 FILLER_98_436 ();
 sg13g2_fill_1 FILLER_98_438 ();
 sg13g2_decap_4 FILLER_98_452 ();
 sg13g2_fill_2 FILLER_98_462 ();
 sg13g2_decap_4 FILLER_98_486 ();
 sg13g2_fill_2 FILLER_98_490 ();
 sg13g2_fill_2 FILLER_98_497 ();
 sg13g2_fill_1 FILLER_98_499 ();
 sg13g2_fill_1 FILLER_98_510 ();
 sg13g2_decap_8 FILLER_98_524 ();
 sg13g2_fill_2 FILLER_98_531 ();
 sg13g2_fill_1 FILLER_98_533 ();
 sg13g2_decap_8 FILLER_98_554 ();
 sg13g2_fill_2 FILLER_98_561 ();
 sg13g2_decap_8 FILLER_98_576 ();
 sg13g2_decap_4 FILLER_98_593 ();
 sg13g2_fill_2 FILLER_98_602 ();
 sg13g2_fill_1 FILLER_98_604 ();
 sg13g2_decap_8 FILLER_98_615 ();
 sg13g2_decap_8 FILLER_98_622 ();
 sg13g2_decap_4 FILLER_98_639 ();
 sg13g2_fill_1 FILLER_98_647 ();
 sg13g2_decap_4 FILLER_98_653 ();
 sg13g2_fill_2 FILLER_98_657 ();
 sg13g2_decap_8 FILLER_98_678 ();
 sg13g2_decap_4 FILLER_98_685 ();
 sg13g2_decap_8 FILLER_98_715 ();
 sg13g2_decap_4 FILLER_98_722 ();
 sg13g2_fill_1 FILLER_98_726 ();
 sg13g2_decap_8 FILLER_98_744 ();
 sg13g2_decap_4 FILLER_98_751 ();
 sg13g2_fill_2 FILLER_98_755 ();
 sg13g2_decap_8 FILLER_98_801 ();
 sg13g2_decap_8 FILLER_98_808 ();
 sg13g2_decap_8 FILLER_98_815 ();
 sg13g2_decap_8 FILLER_98_822 ();
 sg13g2_decap_8 FILLER_98_829 ();
 sg13g2_decap_8 FILLER_98_836 ();
 sg13g2_decap_8 FILLER_98_843 ();
 sg13g2_decap_8 FILLER_98_850 ();
 sg13g2_decap_8 FILLER_98_857 ();
 sg13g2_decap_8 FILLER_98_864 ();
 sg13g2_decap_8 FILLER_98_871 ();
 sg13g2_decap_8 FILLER_98_878 ();
 sg13g2_decap_8 FILLER_98_885 ();
 sg13g2_decap_8 FILLER_98_892 ();
 sg13g2_decap_8 FILLER_98_899 ();
 sg13g2_decap_8 FILLER_98_906 ();
 sg13g2_decap_8 FILLER_98_913 ();
 sg13g2_decap_8 FILLER_98_920 ();
 sg13g2_decap_8 FILLER_98_927 ();
 sg13g2_decap_8 FILLER_98_934 ();
 sg13g2_decap_8 FILLER_98_941 ();
 sg13g2_decap_8 FILLER_98_948 ();
 sg13g2_decap_8 FILLER_98_955 ();
 sg13g2_decap_8 FILLER_98_962 ();
 sg13g2_decap_8 FILLER_98_969 ();
 sg13g2_decap_8 FILLER_98_976 ();
 sg13g2_decap_8 FILLER_98_983 ();
 sg13g2_decap_8 FILLER_98_990 ();
 sg13g2_decap_8 FILLER_98_997 ();
 sg13g2_decap_8 FILLER_98_1004 ();
 sg13g2_decap_8 FILLER_98_1011 ();
 sg13g2_decap_8 FILLER_98_1018 ();
 sg13g2_decap_4 FILLER_98_1025 ();
 sg13g2_decap_8 FILLER_99_0 ();
 sg13g2_decap_8 FILLER_99_7 ();
 sg13g2_decap_8 FILLER_99_14 ();
 sg13g2_decap_8 FILLER_99_21 ();
 sg13g2_decap_8 FILLER_99_28 ();
 sg13g2_decap_8 FILLER_99_35 ();
 sg13g2_decap_8 FILLER_99_42 ();
 sg13g2_decap_8 FILLER_99_49 ();
 sg13g2_decap_8 FILLER_99_56 ();
 sg13g2_decap_8 FILLER_99_63 ();
 sg13g2_decap_8 FILLER_99_70 ();
 sg13g2_decap_8 FILLER_99_77 ();
 sg13g2_decap_8 FILLER_99_84 ();
 sg13g2_decap_8 FILLER_99_91 ();
 sg13g2_decap_8 FILLER_99_98 ();
 sg13g2_decap_8 FILLER_99_105 ();
 sg13g2_decap_8 FILLER_99_112 ();
 sg13g2_decap_8 FILLER_99_119 ();
 sg13g2_decap_8 FILLER_99_126 ();
 sg13g2_decap_8 FILLER_99_133 ();
 sg13g2_decap_8 FILLER_99_140 ();
 sg13g2_decap_4 FILLER_99_147 ();
 sg13g2_fill_2 FILLER_99_160 ();
 sg13g2_decap_8 FILLER_99_171 ();
 sg13g2_decap_8 FILLER_99_178 ();
 sg13g2_fill_1 FILLER_99_194 ();
 sg13g2_decap_8 FILLER_99_232 ();
 sg13g2_fill_2 FILLER_99_239 ();
 sg13g2_fill_1 FILLER_99_241 ();
 sg13g2_decap_8 FILLER_99_252 ();
 sg13g2_fill_1 FILLER_99_259 ();
 sg13g2_fill_1 FILLER_99_269 ();
 sg13g2_decap_8 FILLER_99_280 ();
 sg13g2_fill_1 FILLER_99_287 ();
 sg13g2_decap_8 FILLER_99_297 ();
 sg13g2_decap_8 FILLER_99_304 ();
 sg13g2_fill_1 FILLER_99_311 ();
 sg13g2_fill_1 FILLER_99_341 ();
 sg13g2_decap_8 FILLER_99_351 ();
 sg13g2_decap_8 FILLER_99_358 ();
 sg13g2_decap_8 FILLER_99_365 ();
 sg13g2_decap_8 FILLER_99_372 ();
 sg13g2_decap_8 FILLER_99_379 ();
 sg13g2_decap_8 FILLER_99_386 ();
 sg13g2_fill_2 FILLER_99_393 ();
 sg13g2_fill_1 FILLER_99_395 ();
 sg13g2_decap_8 FILLER_99_417 ();
 sg13g2_decap_8 FILLER_99_424 ();
 sg13g2_fill_2 FILLER_99_431 ();
 sg13g2_fill_1 FILLER_99_433 ();
 sg13g2_fill_2 FILLER_99_442 ();
 sg13g2_fill_1 FILLER_99_444 ();
 sg13g2_decap_8 FILLER_99_463 ();
 sg13g2_fill_1 FILLER_99_470 ();
 sg13g2_decap_8 FILLER_99_490 ();
 sg13g2_fill_2 FILLER_99_497 ();
 sg13g2_decap_4 FILLER_99_503 ();
 sg13g2_decap_4 FILLER_99_528 ();
 sg13g2_fill_2 FILLER_99_532 ();
 sg13g2_fill_2 FILLER_99_538 ();
 sg13g2_fill_1 FILLER_99_540 ();
 sg13g2_decap_4 FILLER_99_552 ();
 sg13g2_fill_1 FILLER_99_556 ();
 sg13g2_decap_4 FILLER_99_562 ();
 sg13g2_fill_1 FILLER_99_566 ();
 sg13g2_fill_2 FILLER_99_572 ();
 sg13g2_fill_2 FILLER_99_629 ();
 sg13g2_fill_2 FILLER_99_644 ();
 sg13g2_fill_1 FILLER_99_657 ();
 sg13g2_decap_8 FILLER_99_681 ();
 sg13g2_decap_8 FILLER_99_688 ();
 sg13g2_fill_1 FILLER_99_695 ();
 sg13g2_decap_8 FILLER_99_712 ();
 sg13g2_decap_8 FILLER_99_719 ();
 sg13g2_fill_2 FILLER_99_726 ();
 sg13g2_fill_2 FILLER_99_743 ();
 sg13g2_decap_4 FILLER_99_762 ();
 sg13g2_decap_8 FILLER_99_790 ();
 sg13g2_decap_8 FILLER_99_797 ();
 sg13g2_decap_8 FILLER_99_804 ();
 sg13g2_decap_8 FILLER_99_811 ();
 sg13g2_decap_8 FILLER_99_818 ();
 sg13g2_decap_8 FILLER_99_825 ();
 sg13g2_decap_8 FILLER_99_832 ();
 sg13g2_decap_8 FILLER_99_839 ();
 sg13g2_decap_8 FILLER_99_846 ();
 sg13g2_decap_8 FILLER_99_853 ();
 sg13g2_decap_8 FILLER_99_860 ();
 sg13g2_decap_8 FILLER_99_867 ();
 sg13g2_decap_8 FILLER_99_874 ();
 sg13g2_decap_8 FILLER_99_881 ();
 sg13g2_decap_8 FILLER_99_888 ();
 sg13g2_decap_8 FILLER_99_895 ();
 sg13g2_decap_8 FILLER_99_902 ();
 sg13g2_decap_8 FILLER_99_909 ();
 sg13g2_decap_8 FILLER_99_916 ();
 sg13g2_decap_8 FILLER_99_923 ();
 sg13g2_decap_8 FILLER_99_930 ();
 sg13g2_decap_8 FILLER_99_937 ();
 sg13g2_decap_8 FILLER_99_944 ();
 sg13g2_decap_8 FILLER_99_951 ();
 sg13g2_decap_8 FILLER_99_958 ();
 sg13g2_decap_8 FILLER_99_965 ();
 sg13g2_decap_8 FILLER_99_972 ();
 sg13g2_decap_8 FILLER_99_979 ();
 sg13g2_decap_8 FILLER_99_986 ();
 sg13g2_decap_8 FILLER_99_993 ();
 sg13g2_decap_8 FILLER_99_1000 ();
 sg13g2_decap_8 FILLER_99_1007 ();
 sg13g2_decap_8 FILLER_99_1014 ();
 sg13g2_decap_8 FILLER_99_1021 ();
 sg13g2_fill_1 FILLER_99_1028 ();
 sg13g2_decap_8 FILLER_100_0 ();
 sg13g2_decap_8 FILLER_100_7 ();
 sg13g2_decap_8 FILLER_100_14 ();
 sg13g2_decap_8 FILLER_100_21 ();
 sg13g2_decap_8 FILLER_100_28 ();
 sg13g2_decap_8 FILLER_100_35 ();
 sg13g2_decap_8 FILLER_100_42 ();
 sg13g2_decap_8 FILLER_100_49 ();
 sg13g2_decap_8 FILLER_100_56 ();
 sg13g2_decap_8 FILLER_100_63 ();
 sg13g2_decap_8 FILLER_100_70 ();
 sg13g2_decap_8 FILLER_100_77 ();
 sg13g2_decap_8 FILLER_100_84 ();
 sg13g2_decap_8 FILLER_100_91 ();
 sg13g2_decap_8 FILLER_100_98 ();
 sg13g2_decap_8 FILLER_100_105 ();
 sg13g2_decap_8 FILLER_100_112 ();
 sg13g2_decap_8 FILLER_100_119 ();
 sg13g2_decap_8 FILLER_100_126 ();
 sg13g2_decap_8 FILLER_100_133 ();
 sg13g2_decap_8 FILLER_100_140 ();
 sg13g2_decap_8 FILLER_100_147 ();
 sg13g2_decap_8 FILLER_100_154 ();
 sg13g2_decap_8 FILLER_100_170 ();
 sg13g2_decap_8 FILLER_100_177 ();
 sg13g2_decap_8 FILLER_100_184 ();
 sg13g2_decap_8 FILLER_100_191 ();
 sg13g2_decap_8 FILLER_100_198 ();
 sg13g2_decap_8 FILLER_100_205 ();
 sg13g2_decap_8 FILLER_100_212 ();
 sg13g2_decap_8 FILLER_100_219 ();
 sg13g2_decap_8 FILLER_100_226 ();
 sg13g2_decap_8 FILLER_100_233 ();
 sg13g2_decap_8 FILLER_100_240 ();
 sg13g2_decap_8 FILLER_100_247 ();
 sg13g2_decap_8 FILLER_100_254 ();
 sg13g2_decap_8 FILLER_100_261 ();
 sg13g2_decap_8 FILLER_100_268 ();
 sg13g2_decap_8 FILLER_100_275 ();
 sg13g2_decap_8 FILLER_100_282 ();
 sg13g2_decap_8 FILLER_100_289 ();
 sg13g2_decap_8 FILLER_100_296 ();
 sg13g2_decap_8 FILLER_100_303 ();
 sg13g2_decap_8 FILLER_100_310 ();
 sg13g2_decap_8 FILLER_100_317 ();
 sg13g2_decap_8 FILLER_100_324 ();
 sg13g2_decap_8 FILLER_100_331 ();
 sg13g2_decap_8 FILLER_100_338 ();
 sg13g2_decap_8 FILLER_100_345 ();
 sg13g2_decap_8 FILLER_100_352 ();
 sg13g2_decap_8 FILLER_100_359 ();
 sg13g2_decap_8 FILLER_100_366 ();
 sg13g2_decap_8 FILLER_100_373 ();
 sg13g2_decap_8 FILLER_100_380 ();
 sg13g2_fill_1 FILLER_100_387 ();
 sg13g2_fill_1 FILLER_100_409 ();
 sg13g2_fill_2 FILLER_100_425 ();
 sg13g2_fill_1 FILLER_100_427 ();
 sg13g2_fill_2 FILLER_100_454 ();
 sg13g2_fill_1 FILLER_100_456 ();
 sg13g2_decap_8 FILLER_100_470 ();
 sg13g2_fill_2 FILLER_100_477 ();
 sg13g2_decap_4 FILLER_100_492 ();
 sg13g2_fill_2 FILLER_100_514 ();
 sg13g2_fill_1 FILLER_100_516 ();
 sg13g2_decap_8 FILLER_100_527 ();
 sg13g2_decap_8 FILLER_100_534 ();
 sg13g2_decap_4 FILLER_100_541 ();
 sg13g2_decap_4 FILLER_100_563 ();
 sg13g2_fill_1 FILLER_100_567 ();
 sg13g2_fill_2 FILLER_100_575 ();
 sg13g2_decap_4 FILLER_100_590 ();
 sg13g2_fill_1 FILLER_100_594 ();
 sg13g2_decap_8 FILLER_100_619 ();
 sg13g2_decap_8 FILLER_100_626 ();
 sg13g2_decap_8 FILLER_100_633 ();
 sg13g2_fill_2 FILLER_100_645 ();
 sg13g2_fill_1 FILLER_100_647 ();
 sg13g2_fill_2 FILLER_100_658 ();
 sg13g2_fill_2 FILLER_100_675 ();
 sg13g2_decap_8 FILLER_100_681 ();
 sg13g2_decap_4 FILLER_100_688 ();
 sg13g2_fill_1 FILLER_100_692 ();
 sg13g2_decap_8 FILLER_100_740 ();
 sg13g2_decap_4 FILLER_100_747 ();
 sg13g2_decap_8 FILLER_100_756 ();
 sg13g2_fill_2 FILLER_100_763 ();
 sg13g2_fill_1 FILLER_100_765 ();
 sg13g2_decap_8 FILLER_100_784 ();
 sg13g2_decap_8 FILLER_100_791 ();
 sg13g2_decap_8 FILLER_100_798 ();
 sg13g2_decap_8 FILLER_100_805 ();
 sg13g2_decap_8 FILLER_100_812 ();
 sg13g2_decap_8 FILLER_100_819 ();
 sg13g2_decap_8 FILLER_100_826 ();
 sg13g2_decap_8 FILLER_100_833 ();
 sg13g2_decap_8 FILLER_100_840 ();
 sg13g2_decap_8 FILLER_100_847 ();
 sg13g2_decap_8 FILLER_100_854 ();
 sg13g2_decap_8 FILLER_100_861 ();
 sg13g2_decap_8 FILLER_100_868 ();
 sg13g2_decap_8 FILLER_100_875 ();
 sg13g2_decap_8 FILLER_100_882 ();
 sg13g2_decap_8 FILLER_100_889 ();
 sg13g2_decap_8 FILLER_100_896 ();
 sg13g2_decap_8 FILLER_100_903 ();
 sg13g2_decap_8 FILLER_100_910 ();
 sg13g2_decap_8 FILLER_100_917 ();
 sg13g2_decap_8 FILLER_100_924 ();
 sg13g2_decap_8 FILLER_100_931 ();
 sg13g2_decap_8 FILLER_100_938 ();
 sg13g2_decap_8 FILLER_100_945 ();
 sg13g2_decap_8 FILLER_100_952 ();
 sg13g2_decap_8 FILLER_100_959 ();
 sg13g2_decap_8 FILLER_100_966 ();
 sg13g2_decap_8 FILLER_100_973 ();
 sg13g2_decap_8 FILLER_100_980 ();
 sg13g2_decap_8 FILLER_100_987 ();
 sg13g2_decap_8 FILLER_100_994 ();
 sg13g2_decap_8 FILLER_100_1001 ();
 sg13g2_decap_8 FILLER_100_1008 ();
 sg13g2_decap_8 FILLER_100_1015 ();
 sg13g2_decap_8 FILLER_100_1022 ();
 sg13g2_decap_8 FILLER_101_0 ();
 sg13g2_decap_8 FILLER_101_7 ();
 sg13g2_decap_8 FILLER_101_14 ();
 sg13g2_decap_8 FILLER_101_21 ();
 sg13g2_decap_8 FILLER_101_28 ();
 sg13g2_decap_8 FILLER_101_35 ();
 sg13g2_decap_8 FILLER_101_42 ();
 sg13g2_decap_8 FILLER_101_49 ();
 sg13g2_decap_8 FILLER_101_56 ();
 sg13g2_decap_8 FILLER_101_63 ();
 sg13g2_decap_8 FILLER_101_70 ();
 sg13g2_decap_8 FILLER_101_77 ();
 sg13g2_decap_8 FILLER_101_84 ();
 sg13g2_decap_8 FILLER_101_91 ();
 sg13g2_decap_8 FILLER_101_98 ();
 sg13g2_decap_8 FILLER_101_105 ();
 sg13g2_decap_8 FILLER_101_112 ();
 sg13g2_decap_8 FILLER_101_119 ();
 sg13g2_decap_8 FILLER_101_126 ();
 sg13g2_decap_8 FILLER_101_133 ();
 sg13g2_decap_8 FILLER_101_140 ();
 sg13g2_decap_8 FILLER_101_147 ();
 sg13g2_decap_8 FILLER_101_154 ();
 sg13g2_decap_8 FILLER_101_161 ();
 sg13g2_decap_8 FILLER_101_168 ();
 sg13g2_decap_8 FILLER_101_175 ();
 sg13g2_decap_8 FILLER_101_182 ();
 sg13g2_decap_8 FILLER_101_189 ();
 sg13g2_decap_8 FILLER_101_196 ();
 sg13g2_decap_8 FILLER_101_203 ();
 sg13g2_decap_8 FILLER_101_210 ();
 sg13g2_decap_8 FILLER_101_217 ();
 sg13g2_decap_8 FILLER_101_224 ();
 sg13g2_decap_8 FILLER_101_231 ();
 sg13g2_decap_8 FILLER_101_238 ();
 sg13g2_decap_8 FILLER_101_245 ();
 sg13g2_decap_8 FILLER_101_252 ();
 sg13g2_decap_8 FILLER_101_259 ();
 sg13g2_decap_8 FILLER_101_266 ();
 sg13g2_decap_8 FILLER_101_273 ();
 sg13g2_decap_8 FILLER_101_280 ();
 sg13g2_decap_8 FILLER_101_287 ();
 sg13g2_decap_8 FILLER_101_294 ();
 sg13g2_decap_8 FILLER_101_301 ();
 sg13g2_decap_8 FILLER_101_308 ();
 sg13g2_decap_8 FILLER_101_315 ();
 sg13g2_decap_8 FILLER_101_322 ();
 sg13g2_decap_8 FILLER_101_329 ();
 sg13g2_decap_8 FILLER_101_336 ();
 sg13g2_decap_8 FILLER_101_343 ();
 sg13g2_decap_8 FILLER_101_350 ();
 sg13g2_decap_8 FILLER_101_357 ();
 sg13g2_decap_8 FILLER_101_364 ();
 sg13g2_decap_8 FILLER_101_371 ();
 sg13g2_decap_8 FILLER_101_378 ();
 sg13g2_decap_4 FILLER_101_385 ();
 sg13g2_fill_1 FILLER_101_389 ();
 sg13g2_decap_8 FILLER_101_425 ();
 sg13g2_decap_8 FILLER_101_432 ();
 sg13g2_fill_2 FILLER_101_459 ();
 sg13g2_decap_4 FILLER_101_471 ();
 sg13g2_fill_2 FILLER_101_475 ();
 sg13g2_fill_2 FILLER_101_492 ();
 sg13g2_fill_1 FILLER_101_503 ();
 sg13g2_fill_2 FILLER_101_518 ();
 sg13g2_fill_1 FILLER_101_520 ();
 sg13g2_fill_1 FILLER_101_529 ();
 sg13g2_decap_8 FILLER_101_534 ();
 sg13g2_decap_4 FILLER_101_541 ();
 sg13g2_fill_1 FILLER_101_545 ();
 sg13g2_fill_2 FILLER_101_562 ();
 sg13g2_fill_1 FILLER_101_564 ();
 sg13g2_fill_2 FILLER_101_578 ();
 sg13g2_fill_1 FILLER_101_580 ();
 sg13g2_decap_4 FILLER_101_585 ();
 sg13g2_fill_1 FILLER_101_589 ();
 sg13g2_fill_2 FILLER_101_595 ();
 sg13g2_decap_4 FILLER_101_601 ();
 sg13g2_decap_8 FILLER_101_609 ();
 sg13g2_fill_2 FILLER_101_633 ();
 sg13g2_fill_1 FILLER_101_640 ();
 sg13g2_fill_1 FILLER_101_656 ();
 sg13g2_fill_1 FILLER_101_662 ();
 sg13g2_decap_4 FILLER_101_668 ();
 sg13g2_fill_1 FILLER_101_672 ();
 sg13g2_fill_2 FILLER_101_683 ();
 sg13g2_fill_1 FILLER_101_685 ();
 sg13g2_decap_8 FILLER_101_691 ();
 sg13g2_decap_4 FILLER_101_698 ();
 sg13g2_fill_2 FILLER_101_702 ();
 sg13g2_decap_8 FILLER_101_708 ();
 sg13g2_decap_8 FILLER_101_715 ();
 sg13g2_decap_4 FILLER_101_722 ();
 sg13g2_fill_1 FILLER_101_726 ();
 sg13g2_decap_8 FILLER_101_746 ();
 sg13g2_decap_4 FILLER_101_753 ();
 sg13g2_fill_2 FILLER_101_761 ();
 sg13g2_decap_8 FILLER_101_791 ();
 sg13g2_decap_8 FILLER_101_798 ();
 sg13g2_decap_8 FILLER_101_805 ();
 sg13g2_decap_8 FILLER_101_812 ();
 sg13g2_decap_8 FILLER_101_819 ();
 sg13g2_decap_8 FILLER_101_826 ();
 sg13g2_decap_8 FILLER_101_833 ();
 sg13g2_decap_8 FILLER_101_840 ();
 sg13g2_decap_8 FILLER_101_847 ();
 sg13g2_decap_8 FILLER_101_854 ();
 sg13g2_decap_8 FILLER_101_861 ();
 sg13g2_decap_8 FILLER_101_868 ();
 sg13g2_decap_8 FILLER_101_875 ();
 sg13g2_decap_8 FILLER_101_882 ();
 sg13g2_decap_8 FILLER_101_889 ();
 sg13g2_decap_8 FILLER_101_896 ();
 sg13g2_decap_8 FILLER_101_903 ();
 sg13g2_decap_8 FILLER_101_910 ();
 sg13g2_decap_8 FILLER_101_917 ();
 sg13g2_decap_8 FILLER_101_924 ();
 sg13g2_decap_8 FILLER_101_931 ();
 sg13g2_decap_8 FILLER_101_938 ();
 sg13g2_decap_8 FILLER_101_945 ();
 sg13g2_decap_8 FILLER_101_952 ();
 sg13g2_decap_8 FILLER_101_959 ();
 sg13g2_decap_8 FILLER_101_966 ();
 sg13g2_decap_8 FILLER_101_973 ();
 sg13g2_decap_8 FILLER_101_980 ();
 sg13g2_decap_8 FILLER_101_987 ();
 sg13g2_decap_8 FILLER_101_994 ();
 sg13g2_decap_8 FILLER_101_1001 ();
 sg13g2_decap_8 FILLER_101_1008 ();
 sg13g2_decap_8 FILLER_101_1015 ();
 sg13g2_decap_8 FILLER_101_1022 ();
 sg13g2_decap_8 FILLER_102_0 ();
 sg13g2_decap_8 FILLER_102_7 ();
 sg13g2_decap_8 FILLER_102_14 ();
 sg13g2_decap_8 FILLER_102_21 ();
 sg13g2_decap_8 FILLER_102_28 ();
 sg13g2_decap_8 FILLER_102_35 ();
 sg13g2_decap_8 FILLER_102_42 ();
 sg13g2_decap_8 FILLER_102_49 ();
 sg13g2_decap_8 FILLER_102_56 ();
 sg13g2_decap_8 FILLER_102_63 ();
 sg13g2_decap_8 FILLER_102_70 ();
 sg13g2_decap_8 FILLER_102_77 ();
 sg13g2_decap_8 FILLER_102_84 ();
 sg13g2_decap_8 FILLER_102_91 ();
 sg13g2_decap_8 FILLER_102_98 ();
 sg13g2_decap_8 FILLER_102_105 ();
 sg13g2_decap_8 FILLER_102_112 ();
 sg13g2_decap_8 FILLER_102_119 ();
 sg13g2_decap_8 FILLER_102_126 ();
 sg13g2_decap_8 FILLER_102_133 ();
 sg13g2_decap_8 FILLER_102_140 ();
 sg13g2_decap_8 FILLER_102_147 ();
 sg13g2_decap_8 FILLER_102_154 ();
 sg13g2_decap_8 FILLER_102_161 ();
 sg13g2_decap_8 FILLER_102_168 ();
 sg13g2_decap_8 FILLER_102_175 ();
 sg13g2_decap_8 FILLER_102_182 ();
 sg13g2_decap_8 FILLER_102_189 ();
 sg13g2_decap_8 FILLER_102_196 ();
 sg13g2_decap_8 FILLER_102_203 ();
 sg13g2_decap_8 FILLER_102_210 ();
 sg13g2_decap_8 FILLER_102_217 ();
 sg13g2_decap_8 FILLER_102_224 ();
 sg13g2_decap_8 FILLER_102_231 ();
 sg13g2_decap_8 FILLER_102_238 ();
 sg13g2_decap_8 FILLER_102_245 ();
 sg13g2_decap_8 FILLER_102_252 ();
 sg13g2_decap_8 FILLER_102_259 ();
 sg13g2_decap_8 FILLER_102_266 ();
 sg13g2_decap_8 FILLER_102_273 ();
 sg13g2_decap_8 FILLER_102_280 ();
 sg13g2_decap_8 FILLER_102_287 ();
 sg13g2_decap_8 FILLER_102_294 ();
 sg13g2_decap_8 FILLER_102_301 ();
 sg13g2_decap_8 FILLER_102_308 ();
 sg13g2_decap_8 FILLER_102_315 ();
 sg13g2_decap_8 FILLER_102_322 ();
 sg13g2_decap_8 FILLER_102_329 ();
 sg13g2_decap_8 FILLER_102_336 ();
 sg13g2_decap_8 FILLER_102_343 ();
 sg13g2_decap_8 FILLER_102_350 ();
 sg13g2_decap_8 FILLER_102_357 ();
 sg13g2_decap_8 FILLER_102_364 ();
 sg13g2_decap_8 FILLER_102_371 ();
 sg13g2_decap_8 FILLER_102_378 ();
 sg13g2_decap_8 FILLER_102_385 ();
 sg13g2_decap_8 FILLER_102_392 ();
 sg13g2_fill_2 FILLER_102_399 ();
 sg13g2_decap_4 FILLER_102_431 ();
 sg13g2_fill_2 FILLER_102_448 ();
 sg13g2_decap_8 FILLER_102_470 ();
 sg13g2_decap_4 FILLER_102_477 ();
 sg13g2_fill_2 FILLER_102_481 ();
 sg13g2_decap_8 FILLER_102_507 ();
 sg13g2_decap_4 FILLER_102_514 ();
 sg13g2_fill_2 FILLER_102_528 ();
 sg13g2_decap_8 FILLER_102_539 ();
 sg13g2_decap_8 FILLER_102_546 ();
 sg13g2_decap_4 FILLER_102_571 ();
 sg13g2_fill_1 FILLER_102_575 ();
 sg13g2_fill_2 FILLER_102_586 ();
 sg13g2_decap_4 FILLER_102_607 ();
 sg13g2_fill_2 FILLER_102_616 ();
 sg13g2_fill_2 FILLER_102_627 ();
 sg13g2_decap_8 FILLER_102_648 ();
 sg13g2_decap_8 FILLER_102_655 ();
 sg13g2_fill_1 FILLER_102_662 ();
 sg13g2_fill_2 FILLER_102_668 ();
 sg13g2_fill_1 FILLER_102_674 ();
 sg13g2_fill_2 FILLER_102_679 ();
 sg13g2_decap_8 FILLER_102_695 ();
 sg13g2_decap_8 FILLER_102_702 ();
 sg13g2_decap_8 FILLER_102_709 ();
 sg13g2_decap_4 FILLER_102_716 ();
 sg13g2_fill_2 FILLER_102_720 ();
 sg13g2_decap_8 FILLER_102_741 ();
 sg13g2_decap_4 FILLER_102_748 ();
 sg13g2_fill_2 FILLER_102_752 ();
 sg13g2_fill_2 FILLER_102_758 ();
 sg13g2_fill_1 FILLER_102_765 ();
 sg13g2_fill_1 FILLER_102_776 ();
 sg13g2_decap_8 FILLER_102_786 ();
 sg13g2_decap_8 FILLER_102_793 ();
 sg13g2_decap_8 FILLER_102_800 ();
 sg13g2_decap_8 FILLER_102_807 ();
 sg13g2_decap_8 FILLER_102_814 ();
 sg13g2_decap_8 FILLER_102_821 ();
 sg13g2_decap_8 FILLER_102_828 ();
 sg13g2_decap_8 FILLER_102_835 ();
 sg13g2_decap_8 FILLER_102_842 ();
 sg13g2_decap_8 FILLER_102_849 ();
 sg13g2_decap_8 FILLER_102_856 ();
 sg13g2_decap_8 FILLER_102_863 ();
 sg13g2_decap_8 FILLER_102_870 ();
 sg13g2_decap_8 FILLER_102_877 ();
 sg13g2_decap_8 FILLER_102_884 ();
 sg13g2_decap_8 FILLER_102_891 ();
 sg13g2_decap_8 FILLER_102_898 ();
 sg13g2_decap_8 FILLER_102_905 ();
 sg13g2_decap_8 FILLER_102_912 ();
 sg13g2_decap_8 FILLER_102_919 ();
 sg13g2_decap_8 FILLER_102_926 ();
 sg13g2_decap_8 FILLER_102_933 ();
 sg13g2_decap_8 FILLER_102_940 ();
 sg13g2_decap_8 FILLER_102_947 ();
 sg13g2_decap_8 FILLER_102_954 ();
 sg13g2_decap_8 FILLER_102_961 ();
 sg13g2_decap_8 FILLER_102_968 ();
 sg13g2_decap_8 FILLER_102_975 ();
 sg13g2_decap_8 FILLER_102_982 ();
 sg13g2_decap_8 FILLER_102_989 ();
 sg13g2_decap_8 FILLER_102_996 ();
 sg13g2_decap_8 FILLER_102_1003 ();
 sg13g2_decap_8 FILLER_102_1010 ();
 sg13g2_decap_8 FILLER_102_1017 ();
 sg13g2_decap_4 FILLER_102_1024 ();
 sg13g2_fill_1 FILLER_102_1028 ();
 sg13g2_decap_8 FILLER_103_0 ();
 sg13g2_decap_8 FILLER_103_7 ();
 sg13g2_decap_8 FILLER_103_14 ();
 sg13g2_decap_8 FILLER_103_21 ();
 sg13g2_decap_8 FILLER_103_28 ();
 sg13g2_decap_8 FILLER_103_35 ();
 sg13g2_decap_8 FILLER_103_42 ();
 sg13g2_decap_8 FILLER_103_49 ();
 sg13g2_decap_8 FILLER_103_56 ();
 sg13g2_decap_8 FILLER_103_63 ();
 sg13g2_decap_8 FILLER_103_70 ();
 sg13g2_decap_8 FILLER_103_77 ();
 sg13g2_decap_8 FILLER_103_84 ();
 sg13g2_decap_8 FILLER_103_91 ();
 sg13g2_decap_8 FILLER_103_98 ();
 sg13g2_decap_8 FILLER_103_105 ();
 sg13g2_decap_8 FILLER_103_112 ();
 sg13g2_decap_8 FILLER_103_119 ();
 sg13g2_decap_8 FILLER_103_126 ();
 sg13g2_decap_8 FILLER_103_133 ();
 sg13g2_decap_8 FILLER_103_140 ();
 sg13g2_decap_8 FILLER_103_147 ();
 sg13g2_decap_8 FILLER_103_154 ();
 sg13g2_decap_8 FILLER_103_161 ();
 sg13g2_decap_8 FILLER_103_168 ();
 sg13g2_decap_8 FILLER_103_175 ();
 sg13g2_decap_8 FILLER_103_182 ();
 sg13g2_decap_8 FILLER_103_189 ();
 sg13g2_decap_8 FILLER_103_196 ();
 sg13g2_decap_8 FILLER_103_203 ();
 sg13g2_decap_8 FILLER_103_210 ();
 sg13g2_decap_8 FILLER_103_217 ();
 sg13g2_decap_8 FILLER_103_224 ();
 sg13g2_decap_8 FILLER_103_231 ();
 sg13g2_decap_8 FILLER_103_238 ();
 sg13g2_decap_8 FILLER_103_245 ();
 sg13g2_decap_8 FILLER_103_252 ();
 sg13g2_decap_8 FILLER_103_259 ();
 sg13g2_decap_8 FILLER_103_266 ();
 sg13g2_decap_8 FILLER_103_273 ();
 sg13g2_decap_8 FILLER_103_280 ();
 sg13g2_decap_8 FILLER_103_287 ();
 sg13g2_decap_8 FILLER_103_294 ();
 sg13g2_decap_8 FILLER_103_301 ();
 sg13g2_decap_8 FILLER_103_308 ();
 sg13g2_decap_8 FILLER_103_315 ();
 sg13g2_decap_8 FILLER_103_322 ();
 sg13g2_decap_8 FILLER_103_329 ();
 sg13g2_decap_8 FILLER_103_336 ();
 sg13g2_decap_8 FILLER_103_343 ();
 sg13g2_decap_8 FILLER_103_350 ();
 sg13g2_decap_8 FILLER_103_357 ();
 sg13g2_decap_8 FILLER_103_364 ();
 sg13g2_decap_8 FILLER_103_371 ();
 sg13g2_decap_8 FILLER_103_378 ();
 sg13g2_decap_8 FILLER_103_385 ();
 sg13g2_decap_8 FILLER_103_392 ();
 sg13g2_decap_8 FILLER_103_399 ();
 sg13g2_decap_8 FILLER_103_406 ();
 sg13g2_fill_2 FILLER_103_413 ();
 sg13g2_fill_1 FILLER_103_415 ();
 sg13g2_decap_8 FILLER_103_421 ();
 sg13g2_fill_1 FILLER_103_428 ();
 sg13g2_fill_1 FILLER_103_472 ();
 sg13g2_fill_1 FILLER_103_481 ();
 sg13g2_fill_1 FILLER_103_486 ();
 sg13g2_fill_2 FILLER_103_496 ();
 sg13g2_fill_1 FILLER_103_498 ();
 sg13g2_decap_4 FILLER_103_504 ();
 sg13g2_fill_1 FILLER_103_508 ();
 sg13g2_fill_2 FILLER_103_518 ();
 sg13g2_fill_1 FILLER_103_520 ();
 sg13g2_fill_1 FILLER_103_525 ();
 sg13g2_decap_8 FILLER_103_530 ();
 sg13g2_fill_1 FILLER_103_537 ();
 sg13g2_fill_2 FILLER_103_542 ();
 sg13g2_fill_1 FILLER_103_544 ();
 sg13g2_fill_2 FILLER_103_550 ();
 sg13g2_decap_8 FILLER_103_557 ();
 sg13g2_decap_8 FILLER_103_564 ();
 sg13g2_decap_8 FILLER_103_571 ();
 sg13g2_fill_2 FILLER_103_603 ();
 sg13g2_decap_4 FILLER_103_618 ();
 sg13g2_fill_1 FILLER_103_622 ();
 sg13g2_fill_1 FILLER_103_629 ();
 sg13g2_fill_1 FILLER_103_639 ();
 sg13g2_decap_8 FILLER_103_644 ();
 sg13g2_decap_4 FILLER_103_651 ();
 sg13g2_fill_1 FILLER_103_655 ();
 sg13g2_fill_2 FILLER_103_671 ();
 sg13g2_decap_8 FILLER_103_701 ();
 sg13g2_decap_8 FILLER_103_708 ();
 sg13g2_fill_2 FILLER_103_715 ();
 sg13g2_decap_4 FILLER_103_737 ();
 sg13g2_fill_2 FILLER_103_751 ();
 sg13g2_fill_1 FILLER_103_762 ();
 sg13g2_fill_2 FILLER_103_767 ();
 sg13g2_fill_1 FILLER_103_769 ();
 sg13g2_decap_8 FILLER_103_774 ();
 sg13g2_decap_8 FILLER_103_781 ();
 sg13g2_decap_8 FILLER_103_788 ();
 sg13g2_decap_8 FILLER_103_795 ();
 sg13g2_decap_8 FILLER_103_802 ();
 sg13g2_decap_8 FILLER_103_809 ();
 sg13g2_decap_8 FILLER_103_816 ();
 sg13g2_decap_8 FILLER_103_823 ();
 sg13g2_decap_8 FILLER_103_830 ();
 sg13g2_decap_8 FILLER_103_837 ();
 sg13g2_decap_8 FILLER_103_844 ();
 sg13g2_decap_8 FILLER_103_851 ();
 sg13g2_decap_8 FILLER_103_858 ();
 sg13g2_decap_8 FILLER_103_865 ();
 sg13g2_decap_8 FILLER_103_872 ();
 sg13g2_decap_8 FILLER_103_879 ();
 sg13g2_decap_8 FILLER_103_886 ();
 sg13g2_decap_8 FILLER_103_893 ();
 sg13g2_decap_8 FILLER_103_900 ();
 sg13g2_decap_8 FILLER_103_907 ();
 sg13g2_decap_8 FILLER_103_914 ();
 sg13g2_decap_8 FILLER_103_921 ();
 sg13g2_decap_8 FILLER_103_928 ();
 sg13g2_decap_8 FILLER_103_935 ();
 sg13g2_decap_8 FILLER_103_942 ();
 sg13g2_decap_8 FILLER_103_949 ();
 sg13g2_decap_8 FILLER_103_956 ();
 sg13g2_decap_8 FILLER_103_963 ();
 sg13g2_decap_8 FILLER_103_970 ();
 sg13g2_decap_8 FILLER_103_977 ();
 sg13g2_decap_8 FILLER_103_984 ();
 sg13g2_decap_8 FILLER_103_991 ();
 sg13g2_decap_8 FILLER_103_998 ();
 sg13g2_decap_8 FILLER_103_1005 ();
 sg13g2_decap_8 FILLER_103_1012 ();
 sg13g2_decap_8 FILLER_103_1019 ();
 sg13g2_fill_2 FILLER_103_1026 ();
 sg13g2_fill_1 FILLER_103_1028 ();
 sg13g2_decap_8 FILLER_104_0 ();
 sg13g2_decap_8 FILLER_104_7 ();
 sg13g2_decap_8 FILLER_104_14 ();
 sg13g2_decap_8 FILLER_104_21 ();
 sg13g2_decap_8 FILLER_104_28 ();
 sg13g2_decap_8 FILLER_104_35 ();
 sg13g2_decap_8 FILLER_104_42 ();
 sg13g2_decap_8 FILLER_104_49 ();
 sg13g2_decap_8 FILLER_104_56 ();
 sg13g2_decap_8 FILLER_104_63 ();
 sg13g2_decap_8 FILLER_104_70 ();
 sg13g2_decap_8 FILLER_104_77 ();
 sg13g2_decap_8 FILLER_104_84 ();
 sg13g2_decap_8 FILLER_104_91 ();
 sg13g2_decap_8 FILLER_104_98 ();
 sg13g2_decap_8 FILLER_104_105 ();
 sg13g2_decap_8 FILLER_104_112 ();
 sg13g2_decap_8 FILLER_104_119 ();
 sg13g2_decap_8 FILLER_104_126 ();
 sg13g2_decap_8 FILLER_104_133 ();
 sg13g2_decap_8 FILLER_104_140 ();
 sg13g2_decap_8 FILLER_104_147 ();
 sg13g2_decap_8 FILLER_104_154 ();
 sg13g2_decap_8 FILLER_104_161 ();
 sg13g2_decap_8 FILLER_104_168 ();
 sg13g2_decap_8 FILLER_104_175 ();
 sg13g2_decap_8 FILLER_104_182 ();
 sg13g2_decap_8 FILLER_104_189 ();
 sg13g2_decap_8 FILLER_104_196 ();
 sg13g2_decap_8 FILLER_104_203 ();
 sg13g2_decap_8 FILLER_104_210 ();
 sg13g2_decap_8 FILLER_104_217 ();
 sg13g2_decap_8 FILLER_104_224 ();
 sg13g2_decap_8 FILLER_104_231 ();
 sg13g2_decap_8 FILLER_104_238 ();
 sg13g2_decap_8 FILLER_104_245 ();
 sg13g2_decap_8 FILLER_104_252 ();
 sg13g2_decap_8 FILLER_104_259 ();
 sg13g2_decap_8 FILLER_104_266 ();
 sg13g2_decap_8 FILLER_104_273 ();
 sg13g2_decap_8 FILLER_104_280 ();
 sg13g2_decap_8 FILLER_104_287 ();
 sg13g2_decap_8 FILLER_104_294 ();
 sg13g2_decap_8 FILLER_104_301 ();
 sg13g2_decap_8 FILLER_104_308 ();
 sg13g2_decap_8 FILLER_104_315 ();
 sg13g2_decap_8 FILLER_104_322 ();
 sg13g2_decap_8 FILLER_104_329 ();
 sg13g2_decap_8 FILLER_104_336 ();
 sg13g2_decap_8 FILLER_104_343 ();
 sg13g2_decap_8 FILLER_104_350 ();
 sg13g2_decap_8 FILLER_104_357 ();
 sg13g2_decap_8 FILLER_104_364 ();
 sg13g2_decap_8 FILLER_104_371 ();
 sg13g2_decap_8 FILLER_104_378 ();
 sg13g2_decap_8 FILLER_104_385 ();
 sg13g2_decap_8 FILLER_104_392 ();
 sg13g2_decap_8 FILLER_104_399 ();
 sg13g2_decap_8 FILLER_104_406 ();
 sg13g2_decap_8 FILLER_104_413 ();
 sg13g2_decap_8 FILLER_104_420 ();
 sg13g2_decap_8 FILLER_104_427 ();
 sg13g2_fill_2 FILLER_104_442 ();
 sg13g2_fill_1 FILLER_104_444 ();
 sg13g2_fill_1 FILLER_104_476 ();
 sg13g2_fill_2 FILLER_104_496 ();
 sg13g2_fill_1 FILLER_104_498 ();
 sg13g2_fill_2 FILLER_104_524 ();
 sg13g2_fill_1 FILLER_104_547 ();
 sg13g2_decap_8 FILLER_104_563 ();
 sg13g2_fill_2 FILLER_104_578 ();
 sg13g2_fill_1 FILLER_104_610 ();
 sg13g2_fill_2 FILLER_104_625 ();
 sg13g2_fill_1 FILLER_104_627 ();
 sg13g2_fill_2 FILLER_104_651 ();
 sg13g2_fill_2 FILLER_104_682 ();
 sg13g2_fill_1 FILLER_104_692 ();
 sg13g2_fill_2 FILLER_104_702 ();
 sg13g2_fill_1 FILLER_104_704 ();
 sg13g2_fill_2 FILLER_104_727 ();
 sg13g2_fill_1 FILLER_104_748 ();
 sg13g2_decap_8 FILLER_104_774 ();
 sg13g2_decap_8 FILLER_104_781 ();
 sg13g2_decap_8 FILLER_104_788 ();
 sg13g2_decap_8 FILLER_104_795 ();
 sg13g2_decap_8 FILLER_104_802 ();
 sg13g2_decap_8 FILLER_104_809 ();
 sg13g2_decap_8 FILLER_104_816 ();
 sg13g2_decap_8 FILLER_104_823 ();
 sg13g2_decap_8 FILLER_104_830 ();
 sg13g2_decap_8 FILLER_104_837 ();
 sg13g2_decap_8 FILLER_104_844 ();
 sg13g2_decap_8 FILLER_104_851 ();
 sg13g2_decap_8 FILLER_104_858 ();
 sg13g2_decap_8 FILLER_104_865 ();
 sg13g2_decap_8 FILLER_104_872 ();
 sg13g2_decap_8 FILLER_104_879 ();
 sg13g2_decap_8 FILLER_104_886 ();
 sg13g2_decap_8 FILLER_104_893 ();
 sg13g2_decap_8 FILLER_104_900 ();
 sg13g2_decap_8 FILLER_104_907 ();
 sg13g2_decap_8 FILLER_104_914 ();
 sg13g2_decap_8 FILLER_104_921 ();
 sg13g2_decap_8 FILLER_104_928 ();
 sg13g2_decap_8 FILLER_104_935 ();
 sg13g2_decap_8 FILLER_104_942 ();
 sg13g2_decap_8 FILLER_104_949 ();
 sg13g2_decap_8 FILLER_104_956 ();
 sg13g2_decap_8 FILLER_104_963 ();
 sg13g2_decap_8 FILLER_104_970 ();
 sg13g2_decap_8 FILLER_104_977 ();
 sg13g2_decap_8 FILLER_104_984 ();
 sg13g2_decap_8 FILLER_104_991 ();
 sg13g2_decap_8 FILLER_104_998 ();
 sg13g2_decap_8 FILLER_104_1005 ();
 sg13g2_decap_8 FILLER_104_1012 ();
 sg13g2_decap_8 FILLER_104_1019 ();
 sg13g2_fill_2 FILLER_104_1026 ();
 sg13g2_fill_1 FILLER_104_1028 ();
 sg13g2_decap_8 FILLER_105_0 ();
 sg13g2_decap_8 FILLER_105_7 ();
 sg13g2_decap_8 FILLER_105_14 ();
 sg13g2_decap_8 FILLER_105_21 ();
 sg13g2_decap_8 FILLER_105_28 ();
 sg13g2_decap_8 FILLER_105_35 ();
 sg13g2_decap_8 FILLER_105_42 ();
 sg13g2_decap_8 FILLER_105_49 ();
 sg13g2_decap_8 FILLER_105_56 ();
 sg13g2_decap_8 FILLER_105_63 ();
 sg13g2_decap_8 FILLER_105_70 ();
 sg13g2_decap_8 FILLER_105_77 ();
 sg13g2_decap_8 FILLER_105_84 ();
 sg13g2_decap_8 FILLER_105_91 ();
 sg13g2_decap_8 FILLER_105_98 ();
 sg13g2_decap_8 FILLER_105_105 ();
 sg13g2_decap_8 FILLER_105_112 ();
 sg13g2_decap_8 FILLER_105_119 ();
 sg13g2_decap_8 FILLER_105_126 ();
 sg13g2_decap_8 FILLER_105_133 ();
 sg13g2_decap_8 FILLER_105_140 ();
 sg13g2_decap_8 FILLER_105_147 ();
 sg13g2_decap_8 FILLER_105_154 ();
 sg13g2_decap_8 FILLER_105_161 ();
 sg13g2_decap_8 FILLER_105_168 ();
 sg13g2_decap_8 FILLER_105_175 ();
 sg13g2_decap_8 FILLER_105_182 ();
 sg13g2_decap_8 FILLER_105_189 ();
 sg13g2_decap_8 FILLER_105_196 ();
 sg13g2_decap_8 FILLER_105_203 ();
 sg13g2_decap_8 FILLER_105_210 ();
 sg13g2_decap_8 FILLER_105_217 ();
 sg13g2_decap_8 FILLER_105_224 ();
 sg13g2_decap_8 FILLER_105_231 ();
 sg13g2_decap_8 FILLER_105_238 ();
 sg13g2_decap_8 FILLER_105_245 ();
 sg13g2_decap_8 FILLER_105_252 ();
 sg13g2_decap_8 FILLER_105_259 ();
 sg13g2_decap_8 FILLER_105_266 ();
 sg13g2_decap_8 FILLER_105_273 ();
 sg13g2_decap_8 FILLER_105_280 ();
 sg13g2_decap_8 FILLER_105_287 ();
 sg13g2_decap_8 FILLER_105_294 ();
 sg13g2_decap_8 FILLER_105_301 ();
 sg13g2_decap_8 FILLER_105_308 ();
 sg13g2_decap_8 FILLER_105_315 ();
 sg13g2_decap_8 FILLER_105_322 ();
 sg13g2_decap_8 FILLER_105_329 ();
 sg13g2_decap_8 FILLER_105_336 ();
 sg13g2_decap_8 FILLER_105_343 ();
 sg13g2_decap_8 FILLER_105_350 ();
 sg13g2_decap_8 FILLER_105_357 ();
 sg13g2_decap_8 FILLER_105_364 ();
 sg13g2_decap_8 FILLER_105_371 ();
 sg13g2_decap_8 FILLER_105_378 ();
 sg13g2_decap_8 FILLER_105_385 ();
 sg13g2_decap_8 FILLER_105_392 ();
 sg13g2_decap_8 FILLER_105_399 ();
 sg13g2_decap_8 FILLER_105_406 ();
 sg13g2_decap_8 FILLER_105_413 ();
 sg13g2_decap_8 FILLER_105_420 ();
 sg13g2_decap_8 FILLER_105_427 ();
 sg13g2_fill_2 FILLER_105_442 ();
 sg13g2_decap_8 FILLER_105_478 ();
 sg13g2_fill_1 FILLER_105_485 ();
 sg13g2_fill_2 FILLER_105_499 ();
 sg13g2_fill_1 FILLER_105_501 ();
 sg13g2_fill_1 FILLER_105_512 ();
 sg13g2_fill_1 FILLER_105_527 ();
 sg13g2_fill_1 FILLER_105_561 ();
 sg13g2_fill_2 FILLER_105_587 ();
 sg13g2_fill_2 FILLER_105_607 ();
 sg13g2_fill_1 FILLER_105_609 ();
 sg13g2_fill_2 FILLER_105_620 ();
 sg13g2_fill_1 FILLER_105_622 ();
 sg13g2_decap_8 FILLER_105_628 ();
 sg13g2_fill_1 FILLER_105_635 ();
 sg13g2_decap_4 FILLER_105_656 ();
 sg13g2_decap_8 FILLER_105_677 ();
 sg13g2_fill_1 FILLER_105_688 ();
 sg13g2_fill_1 FILLER_105_694 ();
 sg13g2_fill_1 FILLER_105_738 ();
 sg13g2_decap_8 FILLER_105_756 ();
 sg13g2_decap_8 FILLER_105_763 ();
 sg13g2_decap_8 FILLER_105_770 ();
 sg13g2_decap_8 FILLER_105_777 ();
 sg13g2_decap_8 FILLER_105_784 ();
 sg13g2_decap_8 FILLER_105_791 ();
 sg13g2_decap_8 FILLER_105_798 ();
 sg13g2_decap_8 FILLER_105_805 ();
 sg13g2_decap_8 FILLER_105_812 ();
 sg13g2_decap_8 FILLER_105_819 ();
 sg13g2_decap_8 FILLER_105_826 ();
 sg13g2_decap_8 FILLER_105_833 ();
 sg13g2_decap_8 FILLER_105_840 ();
 sg13g2_decap_8 FILLER_105_847 ();
 sg13g2_decap_8 FILLER_105_854 ();
 sg13g2_decap_8 FILLER_105_861 ();
 sg13g2_decap_8 FILLER_105_868 ();
 sg13g2_decap_8 FILLER_105_875 ();
 sg13g2_decap_8 FILLER_105_882 ();
 sg13g2_decap_8 FILLER_105_889 ();
 sg13g2_decap_8 FILLER_105_896 ();
 sg13g2_decap_8 FILLER_105_903 ();
 sg13g2_decap_8 FILLER_105_910 ();
 sg13g2_decap_8 FILLER_105_917 ();
 sg13g2_decap_8 FILLER_105_924 ();
 sg13g2_decap_8 FILLER_105_931 ();
 sg13g2_decap_8 FILLER_105_938 ();
 sg13g2_decap_8 FILLER_105_945 ();
 sg13g2_decap_8 FILLER_105_952 ();
 sg13g2_decap_8 FILLER_105_959 ();
 sg13g2_decap_8 FILLER_105_966 ();
 sg13g2_decap_8 FILLER_105_973 ();
 sg13g2_decap_8 FILLER_105_980 ();
 sg13g2_decap_8 FILLER_105_987 ();
 sg13g2_decap_8 FILLER_105_994 ();
 sg13g2_decap_8 FILLER_105_1001 ();
 sg13g2_decap_8 FILLER_105_1008 ();
 sg13g2_decap_8 FILLER_105_1015 ();
 sg13g2_decap_8 FILLER_105_1022 ();
 sg13g2_decap_8 FILLER_106_0 ();
 sg13g2_decap_8 FILLER_106_7 ();
 sg13g2_decap_8 FILLER_106_14 ();
 sg13g2_decap_8 FILLER_106_21 ();
 sg13g2_decap_8 FILLER_106_28 ();
 sg13g2_decap_8 FILLER_106_35 ();
 sg13g2_decap_8 FILLER_106_42 ();
 sg13g2_decap_8 FILLER_106_49 ();
 sg13g2_decap_8 FILLER_106_56 ();
 sg13g2_decap_8 FILLER_106_63 ();
 sg13g2_decap_8 FILLER_106_70 ();
 sg13g2_decap_8 FILLER_106_77 ();
 sg13g2_decap_8 FILLER_106_84 ();
 sg13g2_decap_8 FILLER_106_91 ();
 sg13g2_decap_8 FILLER_106_98 ();
 sg13g2_decap_8 FILLER_106_105 ();
 sg13g2_decap_8 FILLER_106_112 ();
 sg13g2_decap_8 FILLER_106_119 ();
 sg13g2_decap_8 FILLER_106_126 ();
 sg13g2_decap_8 FILLER_106_133 ();
 sg13g2_decap_8 FILLER_106_140 ();
 sg13g2_decap_8 FILLER_106_147 ();
 sg13g2_decap_8 FILLER_106_154 ();
 sg13g2_decap_8 FILLER_106_161 ();
 sg13g2_decap_8 FILLER_106_168 ();
 sg13g2_decap_8 FILLER_106_175 ();
 sg13g2_decap_8 FILLER_106_182 ();
 sg13g2_decap_8 FILLER_106_189 ();
 sg13g2_decap_8 FILLER_106_196 ();
 sg13g2_decap_8 FILLER_106_203 ();
 sg13g2_decap_8 FILLER_106_210 ();
 sg13g2_decap_8 FILLER_106_217 ();
 sg13g2_decap_8 FILLER_106_224 ();
 sg13g2_decap_8 FILLER_106_231 ();
 sg13g2_decap_8 FILLER_106_238 ();
 sg13g2_decap_8 FILLER_106_245 ();
 sg13g2_decap_8 FILLER_106_252 ();
 sg13g2_decap_8 FILLER_106_259 ();
 sg13g2_decap_8 FILLER_106_266 ();
 sg13g2_decap_8 FILLER_106_273 ();
 sg13g2_decap_8 FILLER_106_280 ();
 sg13g2_decap_8 FILLER_106_287 ();
 sg13g2_decap_8 FILLER_106_294 ();
 sg13g2_decap_8 FILLER_106_301 ();
 sg13g2_decap_8 FILLER_106_308 ();
 sg13g2_decap_8 FILLER_106_315 ();
 sg13g2_decap_8 FILLER_106_322 ();
 sg13g2_decap_8 FILLER_106_329 ();
 sg13g2_decap_8 FILLER_106_336 ();
 sg13g2_decap_8 FILLER_106_343 ();
 sg13g2_decap_8 FILLER_106_350 ();
 sg13g2_decap_8 FILLER_106_357 ();
 sg13g2_decap_8 FILLER_106_364 ();
 sg13g2_decap_8 FILLER_106_371 ();
 sg13g2_decap_8 FILLER_106_378 ();
 sg13g2_decap_8 FILLER_106_385 ();
 sg13g2_decap_8 FILLER_106_392 ();
 sg13g2_decap_8 FILLER_106_399 ();
 sg13g2_decap_8 FILLER_106_406 ();
 sg13g2_decap_8 FILLER_106_413 ();
 sg13g2_decap_8 FILLER_106_420 ();
 sg13g2_decap_8 FILLER_106_427 ();
 sg13g2_decap_8 FILLER_106_434 ();
 sg13g2_decap_8 FILLER_106_441 ();
 sg13g2_fill_2 FILLER_106_448 ();
 sg13g2_fill_1 FILLER_106_450 ();
 sg13g2_decap_8 FILLER_106_481 ();
 sg13g2_decap_8 FILLER_106_488 ();
 sg13g2_decap_8 FILLER_106_495 ();
 sg13g2_decap_4 FILLER_106_502 ();
 sg13g2_fill_2 FILLER_106_506 ();
 sg13g2_decap_8 FILLER_106_516 ();
 sg13g2_decap_8 FILLER_106_523 ();
 sg13g2_decap_8 FILLER_106_530 ();
 sg13g2_decap_8 FILLER_106_537 ();
 sg13g2_decap_4 FILLER_106_544 ();
 sg13g2_fill_1 FILLER_106_548 ();
 sg13g2_decap_8 FILLER_106_558 ();
 sg13g2_decap_8 FILLER_106_565 ();
 sg13g2_decap_8 FILLER_106_572 ();
 sg13g2_decap_8 FILLER_106_579 ();
 sg13g2_decap_8 FILLER_106_586 ();
 sg13g2_decap_8 FILLER_106_593 ();
 sg13g2_fill_2 FILLER_106_600 ();
 sg13g2_decap_8 FILLER_106_607 ();
 sg13g2_decap_4 FILLER_106_614 ();
 sg13g2_fill_2 FILLER_106_618 ();
 sg13g2_decap_8 FILLER_106_624 ();
 sg13g2_decap_8 FILLER_106_631 ();
 sg13g2_fill_2 FILLER_106_638 ();
 sg13g2_decap_8 FILLER_106_655 ();
 sg13g2_decap_8 FILLER_106_662 ();
 sg13g2_decap_8 FILLER_106_669 ();
 sg13g2_decap_8 FILLER_106_676 ();
 sg13g2_decap_8 FILLER_106_683 ();
 sg13g2_fill_1 FILLER_106_690 ();
 sg13g2_fill_2 FILLER_106_695 ();
 sg13g2_decap_8 FILLER_106_706 ();
 sg13g2_decap_8 FILLER_106_713 ();
 sg13g2_decap_8 FILLER_106_720 ();
 sg13g2_decap_8 FILLER_106_727 ();
 sg13g2_decap_8 FILLER_106_734 ();
 sg13g2_fill_2 FILLER_106_741 ();
 sg13g2_fill_1 FILLER_106_743 ();
 sg13g2_decap_8 FILLER_106_752 ();
 sg13g2_decap_8 FILLER_106_759 ();
 sg13g2_decap_8 FILLER_106_766 ();
 sg13g2_decap_8 FILLER_106_773 ();
 sg13g2_decap_8 FILLER_106_780 ();
 sg13g2_decap_8 FILLER_106_787 ();
 sg13g2_decap_8 FILLER_106_794 ();
 sg13g2_decap_8 FILLER_106_801 ();
 sg13g2_decap_8 FILLER_106_808 ();
 sg13g2_decap_8 FILLER_106_815 ();
 sg13g2_decap_8 FILLER_106_822 ();
 sg13g2_decap_8 FILLER_106_829 ();
 sg13g2_decap_8 FILLER_106_836 ();
 sg13g2_decap_8 FILLER_106_843 ();
 sg13g2_decap_8 FILLER_106_850 ();
 sg13g2_decap_8 FILLER_106_857 ();
 sg13g2_decap_8 FILLER_106_864 ();
 sg13g2_decap_8 FILLER_106_871 ();
 sg13g2_decap_8 FILLER_106_878 ();
 sg13g2_decap_8 FILLER_106_885 ();
 sg13g2_decap_8 FILLER_106_892 ();
 sg13g2_decap_8 FILLER_106_899 ();
 sg13g2_decap_8 FILLER_106_906 ();
 sg13g2_decap_8 FILLER_106_913 ();
 sg13g2_decap_8 FILLER_106_920 ();
 sg13g2_decap_8 FILLER_106_927 ();
 sg13g2_decap_8 FILLER_106_934 ();
 sg13g2_decap_8 FILLER_106_941 ();
 sg13g2_decap_8 FILLER_106_948 ();
 sg13g2_decap_8 FILLER_106_955 ();
 sg13g2_decap_8 FILLER_106_962 ();
 sg13g2_decap_8 FILLER_106_969 ();
 sg13g2_decap_8 FILLER_106_976 ();
 sg13g2_decap_8 FILLER_106_983 ();
 sg13g2_decap_8 FILLER_106_990 ();
 sg13g2_decap_8 FILLER_106_997 ();
 sg13g2_decap_8 FILLER_106_1004 ();
 sg13g2_decap_8 FILLER_106_1011 ();
 sg13g2_decap_8 FILLER_106_1018 ();
 sg13g2_decap_4 FILLER_106_1025 ();
 assign uio_oe[0] = net32;
 assign uio_oe[1] = net31;
 assign uio_oe[2] = net30;
 assign uio_oe[3] = net29;
 assign uio_oe[4] = net28;
 assign uio_oe[5] = net27;
 assign uio_oe[6] = net26;
 assign uio_oe[7] = net25;
endmodule
