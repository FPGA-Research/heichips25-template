VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO heichips25_snitch_wrapper
  CLASS BLOCK ;
  FOREIGN heichips25_snitch_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 415.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 21.580 3.150 23.780 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 97.180 3.150 99.380 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 172.780 3.150 174.980 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 248.380 3.150 250.580 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 323.980 3.150 326.180 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 399.580 3.150 401.780 408.460 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 475.180 3.150 477.380 408.460 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 15.380 3.560 17.580 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 90.980 3.560 93.180 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 166.580 3.560 168.780 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 242.180 3.560 244.380 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 317.780 3.560 319.980 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 393.380 3.560 395.580 408.870 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 468.980 3.560 471.180 408.870 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 391.660 0.400 392.060 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 382.420 0.400 382.820 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 400.900 0.400 401.300 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.580 0.400 234.980 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 243.820 0.400 244.220 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 253.060 0.400 253.460 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.300 0.400 262.700 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.540 0.400 271.940 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 280.780 0.400 281.180 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 290.020 0.400 290.420 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 299.260 0.400 299.660 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.500 0.400 308.900 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 317.740 0.400 318.140 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.980 0.400 327.380 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.220 0.400 336.620 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 345.460 0.400 345.860 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 354.700 0.400 355.100 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 363.940 0.400 364.340 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 373.180 0.400 373.580 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.660 0.400 161.060 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.900 0.400 170.300 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.140 0.400 179.540 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.380 0.400 188.780 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.620 0.400 198.020 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.860 0.400 207.260 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.100 0.400 216.500 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.340 0.400 225.740 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.400 87.140 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.980 0.400 96.380 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 105.220 0.400 105.620 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.460 0.400 114.860 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.700 0.400 124.100 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.940 0.400 133.340 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.180 0.400 142.580 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.420 0.400 151.820 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.820 0.400 13.220 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.060 0.400 22.460 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.300 0.400 31.700 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.780 0.400 50.180 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.020 0.400 59.420 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 68.260 0.400 68.660 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.500 0.400 77.900 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 496.800 408.390 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 496.800 408.460 ;
      LAYER Metal2 ;
        RECT 0.855 3.635 496.425 408.385 ;
      LAYER Metal3 ;
        RECT 0.400 401.510 496.465 408.340 ;
        RECT 0.610 400.690 496.465 401.510 ;
        RECT 0.400 392.270 496.465 400.690 ;
        RECT 0.610 391.450 496.465 392.270 ;
        RECT 0.400 383.030 496.465 391.450 ;
        RECT 0.610 382.210 496.465 383.030 ;
        RECT 0.400 373.790 496.465 382.210 ;
        RECT 0.610 372.970 496.465 373.790 ;
        RECT 0.400 364.550 496.465 372.970 ;
        RECT 0.610 363.730 496.465 364.550 ;
        RECT 0.400 355.310 496.465 363.730 ;
        RECT 0.610 354.490 496.465 355.310 ;
        RECT 0.400 346.070 496.465 354.490 ;
        RECT 0.610 345.250 496.465 346.070 ;
        RECT 0.400 336.830 496.465 345.250 ;
        RECT 0.610 336.010 496.465 336.830 ;
        RECT 0.400 327.590 496.465 336.010 ;
        RECT 0.610 326.770 496.465 327.590 ;
        RECT 0.400 318.350 496.465 326.770 ;
        RECT 0.610 317.530 496.465 318.350 ;
        RECT 0.400 309.110 496.465 317.530 ;
        RECT 0.610 308.290 496.465 309.110 ;
        RECT 0.400 299.870 496.465 308.290 ;
        RECT 0.610 299.050 496.465 299.870 ;
        RECT 0.400 290.630 496.465 299.050 ;
        RECT 0.610 289.810 496.465 290.630 ;
        RECT 0.400 281.390 496.465 289.810 ;
        RECT 0.610 280.570 496.465 281.390 ;
        RECT 0.400 272.150 496.465 280.570 ;
        RECT 0.610 271.330 496.465 272.150 ;
        RECT 0.400 262.910 496.465 271.330 ;
        RECT 0.610 262.090 496.465 262.910 ;
        RECT 0.400 253.670 496.465 262.090 ;
        RECT 0.610 252.850 496.465 253.670 ;
        RECT 0.400 244.430 496.465 252.850 ;
        RECT 0.610 243.610 496.465 244.430 ;
        RECT 0.400 235.190 496.465 243.610 ;
        RECT 0.610 234.370 496.465 235.190 ;
        RECT 0.400 225.950 496.465 234.370 ;
        RECT 0.610 225.130 496.465 225.950 ;
        RECT 0.400 216.710 496.465 225.130 ;
        RECT 0.610 215.890 496.465 216.710 ;
        RECT 0.400 207.470 496.465 215.890 ;
        RECT 0.610 206.650 496.465 207.470 ;
        RECT 0.400 198.230 496.465 206.650 ;
        RECT 0.610 197.410 496.465 198.230 ;
        RECT 0.400 188.990 496.465 197.410 ;
        RECT 0.610 188.170 496.465 188.990 ;
        RECT 0.400 179.750 496.465 188.170 ;
        RECT 0.610 178.930 496.465 179.750 ;
        RECT 0.400 170.510 496.465 178.930 ;
        RECT 0.610 169.690 496.465 170.510 ;
        RECT 0.400 161.270 496.465 169.690 ;
        RECT 0.610 160.450 496.465 161.270 ;
        RECT 0.400 152.030 496.465 160.450 ;
        RECT 0.610 151.210 496.465 152.030 ;
        RECT 0.400 142.790 496.465 151.210 ;
        RECT 0.610 141.970 496.465 142.790 ;
        RECT 0.400 133.550 496.465 141.970 ;
        RECT 0.610 132.730 496.465 133.550 ;
        RECT 0.400 124.310 496.465 132.730 ;
        RECT 0.610 123.490 496.465 124.310 ;
        RECT 0.400 115.070 496.465 123.490 ;
        RECT 0.610 114.250 496.465 115.070 ;
        RECT 0.400 105.830 496.465 114.250 ;
        RECT 0.610 105.010 496.465 105.830 ;
        RECT 0.400 96.590 496.465 105.010 ;
        RECT 0.610 95.770 496.465 96.590 ;
        RECT 0.400 87.350 496.465 95.770 ;
        RECT 0.610 86.530 496.465 87.350 ;
        RECT 0.400 78.110 496.465 86.530 ;
        RECT 0.610 77.290 496.465 78.110 ;
        RECT 0.400 68.870 496.465 77.290 ;
        RECT 0.610 68.050 496.465 68.870 ;
        RECT 0.400 59.630 496.465 68.050 ;
        RECT 0.610 58.810 496.465 59.630 ;
        RECT 0.400 50.390 496.465 58.810 ;
        RECT 0.610 49.570 496.465 50.390 ;
        RECT 0.400 41.150 496.465 49.570 ;
        RECT 0.610 40.330 496.465 41.150 ;
        RECT 0.400 31.910 496.465 40.330 ;
        RECT 0.610 31.090 496.465 31.910 ;
        RECT 0.400 22.670 496.465 31.090 ;
        RECT 0.610 21.850 496.465 22.670 ;
        RECT 0.400 13.430 496.465 21.850 ;
        RECT 0.610 12.610 496.465 13.430 ;
        RECT 0.400 3.680 496.465 12.610 ;
      LAYER Metal4 ;
        RECT 9.980 3.635 479.140 408.385 ;
      LAYER Metal5 ;
        RECT 15.515 3.470 478.705 408.550 ;
  END
END heichips25_snitch_wrapper
END LIBRARY

