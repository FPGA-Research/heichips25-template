`default_nettype none

module snitch_small_logo ();
endmodule
